magic
tech scmos
timestamp 1554006522
<< ab >>
rect 5 5 45 77
rect 49 5 89 77
rect 93 5 133 77
rect 137 5 177 77
rect 181 5 221 77
rect 225 5 265 77
rect 269 5 309 77
rect 313 5 353 77
rect 357 5 397 77
rect 401 5 441 77
rect 445 5 485 77
rect 489 5 529 77
rect 533 5 573 77
rect 577 5 617 77
rect 621 5 661 77
rect 665 5 705 77
rect 5 -67 408 5
rect 481 -67 666 5
rect 5 -139 659 -67
rect 230 -211 270 -139
rect 274 -211 370 -139
rect 374 -211 470 -139
rect 474 -211 514 -139
rect 518 -211 614 -139
rect 618 -211 714 -139
rect 5 -283 101 -211
rect 105 -283 201 -211
rect 205 -283 245 -211
rect 246 -283 342 -211
rect 346 -283 442 -211
rect 446 -283 486 -211
<< nwell >>
rect 0 37 710 82
rect 0 -62 413 -27
rect 476 -62 671 -27
rect 0 -72 671 -62
rect 0 -107 664 -72
rect 225 -206 719 -171
rect 0 -216 719 -206
rect 0 -251 491 -216
<< pwell >>
rect 0 0 710 37
rect 0 -27 413 0
rect 476 -27 671 0
rect 0 -139 664 -107
rect 0 -144 719 -139
rect 225 -171 719 -144
rect 0 -288 491 -251
<< poly >>
rect 24 62 30 64
rect 24 60 26 62
rect 28 60 30 62
rect 68 62 74 64
rect 68 60 70 62
rect 72 60 74 62
rect 112 62 118 64
rect 112 60 114 62
rect 116 60 118 62
rect 156 62 162 64
rect 156 60 158 62
rect 160 60 162 62
rect 200 62 206 64
rect 200 60 202 62
rect 204 60 206 62
rect 244 62 250 64
rect 244 60 246 62
rect 248 60 250 62
rect 288 62 294 64
rect 288 60 290 62
rect 292 60 294 62
rect 332 62 338 64
rect 332 60 334 62
rect 336 60 338 62
rect 376 62 382 64
rect 376 60 378 62
rect 380 60 382 62
rect 420 62 426 64
rect 420 60 422 62
rect 424 60 426 62
rect 464 62 470 64
rect 464 60 466 62
rect 468 60 470 62
rect 508 62 514 64
rect 508 60 510 62
rect 512 60 514 62
rect 552 62 558 64
rect 552 60 554 62
rect 556 60 558 62
rect 596 62 602 64
rect 596 60 598 62
rect 600 60 602 62
rect 640 62 646 64
rect 640 60 642 62
rect 644 60 646 62
rect 684 62 690 64
rect 684 60 686 62
rect 688 60 690 62
rect 14 55 16 60
rect 24 58 30 60
rect 24 53 26 58
rect 34 53 36 58
rect 58 55 60 60
rect 68 58 74 60
rect 68 53 70 58
rect 78 53 80 58
rect 102 55 104 60
rect 112 58 118 60
rect 112 53 114 58
rect 122 53 124 58
rect 146 55 148 60
rect 156 58 162 60
rect 156 53 158 58
rect 166 53 168 58
rect 190 55 192 60
rect 200 58 206 60
rect 200 53 202 58
rect 210 53 212 58
rect 234 55 236 60
rect 244 58 250 60
rect 244 53 246 58
rect 254 53 256 58
rect 278 55 280 60
rect 288 58 294 60
rect 288 53 290 58
rect 298 53 300 58
rect 322 55 324 60
rect 332 58 338 60
rect 332 53 334 58
rect 342 53 344 58
rect 366 55 368 60
rect 376 58 382 60
rect 376 53 378 58
rect 386 53 388 58
rect 410 55 412 60
rect 420 58 426 60
rect 420 53 422 58
rect 430 53 432 58
rect 454 55 456 60
rect 464 58 470 60
rect 464 53 466 58
rect 474 53 476 58
rect 498 55 500 60
rect 508 58 514 60
rect 508 53 510 58
rect 518 53 520 58
rect 542 55 544 60
rect 552 58 558 60
rect 552 53 554 58
rect 562 53 564 58
rect 586 55 588 60
rect 596 58 602 60
rect 596 53 598 58
rect 606 53 608 58
rect 630 55 632 60
rect 640 58 646 60
rect 640 53 642 58
rect 650 53 652 58
rect 674 55 676 60
rect 684 58 690 60
rect 684 53 686 58
rect 694 53 696 58
rect 14 40 16 43
rect 24 40 26 43
rect 14 38 20 40
rect 14 36 16 38
rect 18 36 20 38
rect 24 37 28 40
rect 14 34 20 36
rect 14 26 16 34
rect 26 23 28 37
rect 34 32 36 43
rect 58 40 60 43
rect 68 40 70 43
rect 58 38 64 40
rect 58 36 60 38
rect 62 36 64 38
rect 68 37 72 40
rect 58 34 64 36
rect 33 30 39 32
rect 33 28 35 30
rect 37 28 39 30
rect 33 26 39 28
rect 58 26 60 34
rect 33 23 35 26
rect 14 16 16 20
rect 70 23 72 37
rect 78 32 80 43
rect 102 40 104 43
rect 112 40 114 43
rect 102 38 108 40
rect 102 36 104 38
rect 106 36 108 38
rect 112 37 116 40
rect 102 34 108 36
rect 77 30 83 32
rect 77 28 79 30
rect 81 28 83 30
rect 77 26 83 28
rect 102 26 104 34
rect 77 23 79 26
rect 58 16 60 20
rect 114 23 116 37
rect 122 32 124 43
rect 146 40 148 43
rect 156 40 158 43
rect 146 38 152 40
rect 146 36 148 38
rect 150 36 152 38
rect 156 37 160 40
rect 146 34 152 36
rect 121 30 127 32
rect 121 28 123 30
rect 125 28 127 30
rect 121 26 127 28
rect 146 26 148 34
rect 121 23 123 26
rect 102 16 104 20
rect 158 23 160 37
rect 166 32 168 43
rect 190 40 192 43
rect 200 40 202 43
rect 190 38 196 40
rect 190 36 192 38
rect 194 36 196 38
rect 200 37 204 40
rect 190 34 196 36
rect 165 30 171 32
rect 165 28 167 30
rect 169 28 171 30
rect 165 26 171 28
rect 190 26 192 34
rect 165 23 167 26
rect 146 16 148 20
rect 202 23 204 37
rect 210 32 212 43
rect 234 40 236 43
rect 244 40 246 43
rect 234 38 240 40
rect 234 36 236 38
rect 238 36 240 38
rect 244 37 248 40
rect 234 34 240 36
rect 209 30 215 32
rect 209 28 211 30
rect 213 28 215 30
rect 209 26 215 28
rect 234 26 236 34
rect 209 23 211 26
rect 190 16 192 20
rect 246 23 248 37
rect 254 32 256 43
rect 278 40 280 43
rect 288 40 290 43
rect 278 38 284 40
rect 278 36 280 38
rect 282 36 284 38
rect 288 37 292 40
rect 278 34 284 36
rect 253 30 259 32
rect 253 28 255 30
rect 257 28 259 30
rect 253 26 259 28
rect 278 26 280 34
rect 253 23 255 26
rect 234 16 236 20
rect 290 23 292 37
rect 298 32 300 43
rect 322 40 324 43
rect 332 40 334 43
rect 322 38 328 40
rect 322 36 324 38
rect 326 36 328 38
rect 332 37 336 40
rect 322 34 328 36
rect 297 30 303 32
rect 297 28 299 30
rect 301 28 303 30
rect 297 26 303 28
rect 322 26 324 34
rect 297 23 299 26
rect 278 16 280 20
rect 334 23 336 37
rect 342 32 344 43
rect 366 40 368 43
rect 376 40 378 43
rect 366 38 372 40
rect 366 36 368 38
rect 370 36 372 38
rect 376 37 380 40
rect 366 34 372 36
rect 341 30 347 32
rect 341 28 343 30
rect 345 28 347 30
rect 341 26 347 28
rect 366 26 368 34
rect 341 23 343 26
rect 322 16 324 20
rect 378 23 380 37
rect 386 32 388 43
rect 410 40 412 43
rect 420 40 422 43
rect 410 38 416 40
rect 410 36 412 38
rect 414 36 416 38
rect 420 37 424 40
rect 410 34 416 36
rect 385 30 391 32
rect 385 28 387 30
rect 389 28 391 30
rect 385 26 391 28
rect 410 26 412 34
rect 385 23 387 26
rect 366 16 368 20
rect 422 23 424 37
rect 430 32 432 43
rect 454 40 456 43
rect 464 40 466 43
rect 454 38 460 40
rect 454 36 456 38
rect 458 36 460 38
rect 464 37 468 40
rect 454 34 460 36
rect 429 30 435 32
rect 429 28 431 30
rect 433 28 435 30
rect 429 26 435 28
rect 454 26 456 34
rect 429 23 431 26
rect 410 16 412 20
rect 466 23 468 37
rect 474 32 476 43
rect 498 40 500 43
rect 508 40 510 43
rect 498 38 504 40
rect 498 36 500 38
rect 502 36 504 38
rect 508 37 512 40
rect 498 34 504 36
rect 473 30 479 32
rect 473 28 475 30
rect 477 28 479 30
rect 473 26 479 28
rect 498 26 500 34
rect 473 23 475 26
rect 454 16 456 20
rect 510 23 512 37
rect 518 32 520 43
rect 542 40 544 43
rect 552 40 554 43
rect 542 38 548 40
rect 542 36 544 38
rect 546 36 548 38
rect 552 37 556 40
rect 542 34 548 36
rect 517 30 523 32
rect 517 28 519 30
rect 521 28 523 30
rect 517 26 523 28
rect 542 26 544 34
rect 517 23 519 26
rect 498 16 500 20
rect 554 23 556 37
rect 562 32 564 43
rect 586 40 588 43
rect 596 40 598 43
rect 586 38 592 40
rect 586 36 588 38
rect 590 36 592 38
rect 596 37 600 40
rect 586 34 592 36
rect 561 30 567 32
rect 561 28 563 30
rect 565 28 567 30
rect 561 26 567 28
rect 586 26 588 34
rect 561 23 563 26
rect 542 16 544 20
rect 598 23 600 37
rect 606 32 608 43
rect 630 40 632 43
rect 640 40 642 43
rect 630 38 636 40
rect 630 36 632 38
rect 634 36 636 38
rect 640 37 644 40
rect 630 34 636 36
rect 605 30 611 32
rect 605 28 607 30
rect 609 28 611 30
rect 605 26 611 28
rect 630 26 632 34
rect 605 23 607 26
rect 586 16 588 20
rect 642 23 644 37
rect 650 32 652 43
rect 674 40 676 43
rect 684 40 686 43
rect 674 38 680 40
rect 674 36 676 38
rect 678 36 680 38
rect 684 37 688 40
rect 674 34 680 36
rect 649 30 655 32
rect 649 28 651 30
rect 653 28 655 30
rect 649 26 655 28
rect 674 26 676 34
rect 649 23 651 26
rect 630 16 632 20
rect 686 23 688 37
rect 694 32 696 43
rect 693 30 699 32
rect 693 28 695 30
rect 697 28 699 30
rect 693 26 699 28
rect 693 23 695 26
rect 674 16 676 20
rect 26 9 28 14
rect 33 9 35 14
rect 70 9 72 14
rect 77 9 79 14
rect 114 9 116 14
rect 121 9 123 14
rect 158 9 160 14
rect 165 9 167 14
rect 202 9 204 14
rect 209 9 211 14
rect 246 9 248 14
rect 253 9 255 14
rect 290 9 292 14
rect 297 9 299 14
rect 334 9 336 14
rect 341 9 343 14
rect 378 9 380 14
rect 385 9 387 14
rect 422 9 424 14
rect 429 9 431 14
rect 466 9 468 14
rect 473 9 475 14
rect 510 9 512 14
rect 517 9 519 14
rect 554 9 556 14
rect 561 9 563 14
rect 598 9 600 14
rect 605 9 607 14
rect 642 9 644 14
rect 649 9 651 14
rect 686 9 688 14
rect 693 9 695 14
rect 22 -1 24 3
rect 33 -1 35 3
rect 40 -1 42 3
rect 22 -24 24 -15
rect 60 -7 62 -2
rect 70 -7 72 -2
rect 80 -4 82 1
rect 90 -1 92 3
rect 111 -1 113 3
rect 122 -1 124 3
rect 129 -1 131 3
rect 33 -24 35 -21
rect 40 -24 42 -21
rect 60 -24 62 -21
rect 70 -24 72 -21
rect 20 -26 26 -24
rect 20 -28 22 -26
rect 24 -28 26 -26
rect 20 -30 26 -28
rect 30 -26 36 -24
rect 30 -28 32 -26
rect 34 -28 36 -26
rect 30 -30 36 -28
rect 40 -26 62 -24
rect 40 -28 42 -26
rect 44 -28 49 -26
rect 51 -28 62 -26
rect 40 -30 62 -28
rect 66 -26 72 -24
rect 66 -28 68 -26
rect 70 -28 72 -26
rect 66 -30 72 -28
rect 80 -27 82 -14
rect 90 -17 92 -14
rect 86 -19 92 -17
rect 86 -21 88 -19
rect 90 -21 92 -19
rect 86 -23 92 -21
rect 80 -29 86 -27
rect 22 -33 24 -30
rect 32 -33 34 -30
rect 42 -33 44 -30
rect 60 -33 62 -30
rect 67 -33 69 -30
rect 80 -31 82 -29
rect 84 -31 86 -29
rect 77 -33 86 -31
rect 77 -36 79 -33
rect 90 -36 92 -23
rect 111 -24 113 -15
rect 149 -7 151 -2
rect 159 -7 161 -2
rect 169 -4 171 1
rect 179 -1 181 3
rect 240 -1 242 3
rect 251 -1 253 3
rect 258 -1 260 3
rect 199 -10 201 -6
rect 209 -10 211 -6
rect 219 -10 221 -6
rect 122 -24 124 -21
rect 129 -24 131 -21
rect 149 -24 151 -21
rect 159 -24 161 -21
rect 109 -26 115 -24
rect 109 -28 111 -26
rect 113 -28 115 -26
rect 109 -30 115 -28
rect 119 -26 125 -24
rect 119 -28 121 -26
rect 123 -28 125 -26
rect 119 -30 125 -28
rect 129 -26 151 -24
rect 129 -28 131 -26
rect 133 -28 138 -26
rect 140 -28 151 -26
rect 129 -30 151 -28
rect 155 -26 161 -24
rect 155 -28 157 -26
rect 159 -28 161 -26
rect 155 -30 161 -28
rect 169 -27 171 -14
rect 179 -17 181 -14
rect 175 -19 181 -17
rect 175 -21 177 -19
rect 179 -21 181 -19
rect 175 -23 181 -21
rect 169 -29 175 -27
rect 111 -33 113 -30
rect 121 -33 123 -30
rect 131 -33 133 -30
rect 149 -33 151 -30
rect 156 -33 158 -30
rect 169 -31 171 -29
rect 173 -31 175 -29
rect 166 -33 175 -31
rect 77 -54 79 -49
rect 22 -65 24 -61
rect 32 -65 34 -61
rect 42 -65 44 -61
rect 60 -63 62 -58
rect 67 -63 69 -58
rect 166 -36 168 -33
rect 179 -36 181 -23
rect 199 -24 201 -16
rect 195 -26 201 -24
rect 195 -28 197 -26
rect 199 -28 201 -26
rect 195 -30 201 -28
rect 166 -54 168 -49
rect 90 -65 92 -61
rect 111 -65 113 -61
rect 121 -65 123 -61
rect 131 -65 133 -61
rect 149 -63 151 -58
rect 156 -63 158 -58
rect 199 -43 201 -30
rect 209 -32 211 -16
rect 219 -25 221 -16
rect 240 -24 242 -15
rect 278 -7 280 -2
rect 288 -7 290 -2
rect 298 -4 300 1
rect 308 -1 310 3
rect 329 -1 331 3
rect 340 -1 342 3
rect 347 -1 349 3
rect 251 -24 253 -21
rect 258 -24 260 -21
rect 278 -24 280 -21
rect 288 -24 290 -21
rect 215 -27 221 -25
rect 215 -29 217 -27
rect 219 -29 221 -27
rect 215 -31 221 -29
rect 238 -26 244 -24
rect 238 -28 240 -26
rect 242 -28 244 -26
rect 238 -30 244 -28
rect 248 -26 254 -24
rect 248 -28 250 -26
rect 252 -28 254 -26
rect 248 -30 254 -28
rect 258 -26 280 -24
rect 258 -28 260 -26
rect 262 -28 267 -26
rect 269 -28 280 -26
rect 258 -30 280 -28
rect 284 -26 290 -24
rect 284 -28 286 -26
rect 288 -28 290 -26
rect 284 -30 290 -28
rect 298 -27 300 -14
rect 308 -17 310 -14
rect 304 -19 310 -17
rect 304 -21 306 -19
rect 308 -21 310 -19
rect 304 -23 310 -21
rect 298 -29 304 -27
rect 205 -34 211 -32
rect 205 -36 207 -34
rect 209 -36 211 -34
rect 205 -38 211 -36
rect 206 -43 208 -38
rect 219 -40 221 -31
rect 240 -33 242 -30
rect 250 -33 252 -30
rect 260 -33 262 -30
rect 278 -33 280 -30
rect 285 -33 287 -30
rect 298 -31 300 -29
rect 302 -31 304 -29
rect 295 -33 304 -31
rect 219 -56 221 -52
rect 179 -65 181 -61
rect 199 -65 201 -61
rect 206 -65 208 -61
rect 295 -36 297 -33
rect 308 -36 310 -23
rect 329 -24 331 -15
rect 367 -7 369 -2
rect 377 -7 379 -2
rect 387 -4 389 1
rect 397 -1 399 3
rect 498 -1 500 3
rect 509 -1 511 3
rect 516 -1 518 3
rect 340 -24 342 -21
rect 347 -24 349 -21
rect 367 -24 369 -21
rect 377 -24 379 -21
rect 327 -26 333 -24
rect 327 -28 329 -26
rect 331 -28 333 -26
rect 327 -30 333 -28
rect 337 -26 343 -24
rect 337 -28 339 -26
rect 341 -28 343 -26
rect 337 -30 343 -28
rect 347 -26 369 -24
rect 347 -28 349 -26
rect 351 -28 356 -26
rect 358 -28 369 -26
rect 347 -30 369 -28
rect 373 -26 379 -24
rect 373 -28 375 -26
rect 377 -28 379 -26
rect 373 -30 379 -28
rect 387 -27 389 -14
rect 397 -17 399 -14
rect 393 -19 399 -17
rect 393 -21 395 -19
rect 397 -21 399 -19
rect 393 -23 399 -21
rect 387 -29 393 -27
rect 329 -33 331 -30
rect 339 -33 341 -30
rect 349 -33 351 -30
rect 367 -33 369 -30
rect 374 -33 376 -30
rect 387 -31 389 -29
rect 391 -31 393 -29
rect 384 -33 393 -31
rect 295 -54 297 -49
rect 240 -65 242 -61
rect 250 -65 252 -61
rect 260 -65 262 -61
rect 278 -63 280 -58
rect 285 -63 287 -58
rect 384 -36 386 -33
rect 397 -36 399 -23
rect 498 -24 500 -15
rect 536 -7 538 -2
rect 546 -7 548 -2
rect 556 -4 558 1
rect 566 -1 568 3
rect 587 -1 589 3
rect 598 -1 600 3
rect 605 -1 607 3
rect 509 -24 511 -21
rect 516 -24 518 -21
rect 536 -24 538 -21
rect 546 -24 548 -21
rect 496 -26 502 -24
rect 496 -28 498 -26
rect 500 -28 502 -26
rect 496 -30 502 -28
rect 506 -26 512 -24
rect 506 -28 508 -26
rect 510 -28 512 -26
rect 506 -30 512 -28
rect 516 -26 538 -24
rect 516 -28 518 -26
rect 520 -28 525 -26
rect 527 -28 538 -26
rect 516 -30 538 -28
rect 542 -26 548 -24
rect 542 -28 544 -26
rect 546 -28 548 -26
rect 542 -30 548 -28
rect 556 -27 558 -14
rect 566 -17 568 -14
rect 562 -19 568 -17
rect 562 -21 564 -19
rect 566 -21 568 -19
rect 562 -23 568 -21
rect 556 -29 562 -27
rect 498 -33 500 -30
rect 508 -33 510 -30
rect 518 -33 520 -30
rect 536 -33 538 -30
rect 543 -33 545 -30
rect 556 -31 558 -29
rect 560 -31 562 -29
rect 553 -33 562 -31
rect 384 -54 386 -49
rect 308 -65 310 -61
rect 329 -65 331 -61
rect 339 -65 341 -61
rect 349 -65 351 -61
rect 367 -63 369 -58
rect 374 -63 376 -58
rect 553 -36 555 -33
rect 566 -36 568 -23
rect 587 -24 589 -15
rect 625 -7 627 -2
rect 635 -7 637 -2
rect 645 -4 647 1
rect 655 -1 657 3
rect 598 -24 600 -21
rect 605 -24 607 -21
rect 625 -24 627 -21
rect 635 -24 637 -21
rect 585 -26 591 -24
rect 585 -28 587 -26
rect 589 -28 591 -26
rect 585 -30 591 -28
rect 595 -26 601 -24
rect 595 -28 597 -26
rect 599 -28 601 -26
rect 595 -30 601 -28
rect 605 -26 627 -24
rect 605 -28 607 -26
rect 609 -28 614 -26
rect 616 -28 627 -26
rect 605 -30 627 -28
rect 631 -26 637 -24
rect 631 -28 633 -26
rect 635 -28 637 -26
rect 631 -30 637 -28
rect 645 -27 647 -14
rect 655 -17 657 -14
rect 651 -19 657 -17
rect 651 -21 653 -19
rect 655 -21 657 -19
rect 651 -23 657 -21
rect 645 -29 651 -27
rect 587 -33 589 -30
rect 597 -33 599 -30
rect 607 -33 609 -30
rect 625 -33 627 -30
rect 632 -33 634 -30
rect 645 -31 647 -29
rect 649 -31 651 -29
rect 642 -33 651 -31
rect 553 -54 555 -49
rect 397 -65 399 -61
rect 498 -65 500 -61
rect 508 -65 510 -61
rect 518 -65 520 -61
rect 536 -63 538 -58
rect 543 -63 545 -58
rect 642 -36 644 -33
rect 655 -36 657 -23
rect 642 -54 644 -49
rect 566 -65 568 -61
rect 587 -65 589 -61
rect 597 -65 599 -61
rect 607 -65 609 -61
rect 625 -63 627 -58
rect 632 -63 634 -58
rect 655 -65 657 -61
rect 14 -73 16 -69
rect 37 -76 39 -71
rect 44 -76 46 -71
rect 62 -73 64 -69
rect 72 -73 74 -69
rect 82 -73 84 -69
rect 103 -73 105 -69
rect 27 -85 29 -80
rect 14 -111 16 -98
rect 27 -101 29 -98
rect 126 -76 128 -71
rect 133 -76 135 -71
rect 151 -73 153 -69
rect 161 -73 163 -69
rect 171 -73 173 -69
rect 116 -85 118 -80
rect 20 -103 29 -101
rect 20 -105 22 -103
rect 24 -105 26 -103
rect 37 -104 39 -101
rect 44 -104 46 -101
rect 62 -104 64 -101
rect 72 -104 74 -101
rect 82 -104 84 -101
rect 20 -107 26 -105
rect 14 -113 20 -111
rect 14 -115 16 -113
rect 18 -115 20 -113
rect 14 -117 20 -115
rect 14 -120 16 -117
rect 24 -120 26 -107
rect 34 -106 40 -104
rect 34 -108 36 -106
rect 38 -108 40 -106
rect 34 -110 40 -108
rect 44 -106 66 -104
rect 44 -108 55 -106
rect 57 -108 62 -106
rect 64 -108 66 -106
rect 44 -110 66 -108
rect 70 -106 76 -104
rect 70 -108 72 -106
rect 74 -108 76 -106
rect 70 -110 76 -108
rect 80 -106 86 -104
rect 80 -108 82 -106
rect 84 -108 86 -106
rect 80 -110 86 -108
rect 34 -113 36 -110
rect 44 -113 46 -110
rect 64 -113 66 -110
rect 71 -113 73 -110
rect 14 -137 16 -133
rect 24 -135 26 -130
rect 34 -132 36 -127
rect 44 -132 46 -127
rect 82 -119 84 -110
rect 103 -111 105 -98
rect 116 -101 118 -98
rect 205 -73 207 -69
rect 212 -73 214 -69
rect 232 -73 234 -69
rect 192 -82 194 -78
rect 109 -103 118 -101
rect 109 -105 111 -103
rect 113 -105 115 -103
rect 126 -104 128 -101
rect 133 -104 135 -101
rect 151 -104 153 -101
rect 161 -104 163 -101
rect 171 -104 173 -101
rect 192 -103 194 -94
rect 205 -96 207 -91
rect 202 -98 208 -96
rect 202 -100 204 -98
rect 206 -100 208 -98
rect 202 -102 208 -100
rect 109 -107 115 -105
rect 103 -113 109 -111
rect 103 -115 105 -113
rect 107 -115 109 -113
rect 103 -117 109 -115
rect 103 -120 105 -117
rect 113 -120 115 -107
rect 123 -106 129 -104
rect 123 -108 125 -106
rect 127 -108 129 -106
rect 123 -110 129 -108
rect 133 -106 155 -104
rect 133 -108 144 -106
rect 146 -108 151 -106
rect 153 -108 155 -106
rect 133 -110 155 -108
rect 159 -106 165 -104
rect 159 -108 161 -106
rect 163 -108 165 -106
rect 159 -110 165 -108
rect 169 -106 175 -104
rect 169 -108 171 -106
rect 173 -108 175 -106
rect 169 -110 175 -108
rect 192 -105 198 -103
rect 192 -107 194 -105
rect 196 -107 198 -105
rect 192 -109 198 -107
rect 123 -113 125 -110
rect 133 -113 135 -110
rect 153 -113 155 -110
rect 160 -113 162 -110
rect 64 -137 66 -133
rect 71 -137 73 -133
rect 82 -137 84 -133
rect 103 -137 105 -133
rect 113 -135 115 -130
rect 123 -132 125 -127
rect 133 -132 135 -127
rect 171 -119 173 -110
rect 192 -118 194 -109
rect 202 -118 204 -102
rect 212 -104 214 -91
rect 255 -76 257 -71
rect 262 -76 264 -71
rect 280 -73 282 -69
rect 290 -73 292 -69
rect 300 -73 302 -69
rect 321 -73 323 -69
rect 245 -85 247 -80
rect 212 -106 218 -104
rect 212 -108 214 -106
rect 216 -108 218 -106
rect 212 -110 218 -108
rect 212 -118 214 -110
rect 232 -111 234 -98
rect 245 -101 247 -98
rect 344 -76 346 -71
rect 351 -76 353 -71
rect 369 -73 371 -69
rect 379 -73 381 -69
rect 389 -73 391 -69
rect 334 -85 336 -80
rect 238 -103 247 -101
rect 238 -105 240 -103
rect 242 -105 244 -103
rect 255 -104 257 -101
rect 262 -104 264 -101
rect 280 -104 282 -101
rect 290 -104 292 -101
rect 300 -104 302 -101
rect 238 -107 244 -105
rect 232 -113 238 -111
rect 232 -115 234 -113
rect 236 -115 238 -113
rect 232 -117 238 -115
rect 232 -120 234 -117
rect 242 -120 244 -107
rect 252 -106 258 -104
rect 252 -108 254 -106
rect 256 -108 258 -106
rect 252 -110 258 -108
rect 262 -106 284 -104
rect 262 -108 273 -106
rect 275 -108 280 -106
rect 282 -108 284 -106
rect 262 -110 284 -108
rect 288 -106 294 -104
rect 288 -108 290 -106
rect 292 -108 294 -106
rect 288 -110 294 -108
rect 298 -106 304 -104
rect 298 -108 300 -106
rect 302 -108 304 -106
rect 298 -110 304 -108
rect 252 -113 254 -110
rect 262 -113 264 -110
rect 282 -113 284 -110
rect 289 -113 291 -110
rect 192 -128 194 -124
rect 202 -128 204 -124
rect 212 -128 214 -124
rect 153 -137 155 -133
rect 160 -137 162 -133
rect 171 -137 173 -133
rect 232 -137 234 -133
rect 242 -135 244 -130
rect 252 -132 254 -127
rect 262 -132 264 -127
rect 300 -119 302 -110
rect 321 -111 323 -98
rect 334 -101 336 -98
rect 423 -73 425 -69
rect 430 -73 432 -69
rect 450 -73 452 -69
rect 410 -82 412 -78
rect 327 -103 336 -101
rect 327 -105 329 -103
rect 331 -105 333 -103
rect 344 -104 346 -101
rect 351 -104 353 -101
rect 369 -104 371 -101
rect 379 -104 381 -101
rect 389 -104 391 -101
rect 410 -103 412 -94
rect 423 -96 425 -91
rect 420 -98 426 -96
rect 420 -100 422 -98
rect 424 -100 426 -98
rect 420 -102 426 -100
rect 327 -107 333 -105
rect 321 -113 327 -111
rect 321 -115 323 -113
rect 325 -115 327 -113
rect 321 -117 327 -115
rect 321 -120 323 -117
rect 331 -120 333 -107
rect 341 -106 347 -104
rect 341 -108 343 -106
rect 345 -108 347 -106
rect 341 -110 347 -108
rect 351 -106 373 -104
rect 351 -108 362 -106
rect 364 -108 369 -106
rect 371 -108 373 -106
rect 351 -110 373 -108
rect 377 -106 383 -104
rect 377 -108 379 -106
rect 381 -108 383 -106
rect 377 -110 383 -108
rect 387 -106 393 -104
rect 387 -108 389 -106
rect 391 -108 393 -106
rect 387 -110 393 -108
rect 410 -105 416 -103
rect 410 -107 412 -105
rect 414 -107 416 -105
rect 410 -109 416 -107
rect 341 -113 343 -110
rect 351 -113 353 -110
rect 371 -113 373 -110
rect 378 -113 380 -110
rect 282 -137 284 -133
rect 289 -137 291 -133
rect 300 -137 302 -133
rect 321 -137 323 -133
rect 331 -135 333 -130
rect 341 -132 343 -127
rect 351 -132 353 -127
rect 389 -119 391 -110
rect 410 -118 412 -109
rect 420 -118 422 -102
rect 430 -104 432 -91
rect 473 -76 475 -71
rect 480 -76 482 -71
rect 498 -73 500 -69
rect 508 -73 510 -69
rect 518 -73 520 -69
rect 539 -73 541 -69
rect 463 -85 465 -80
rect 430 -106 436 -104
rect 430 -108 432 -106
rect 434 -108 436 -106
rect 430 -110 436 -108
rect 430 -118 432 -110
rect 450 -111 452 -98
rect 463 -101 465 -98
rect 562 -76 564 -71
rect 569 -76 571 -71
rect 587 -73 589 -69
rect 597 -73 599 -69
rect 607 -73 609 -69
rect 552 -85 554 -80
rect 456 -103 465 -101
rect 456 -105 458 -103
rect 460 -105 462 -103
rect 473 -104 475 -101
rect 480 -104 482 -101
rect 498 -104 500 -101
rect 508 -104 510 -101
rect 518 -104 520 -101
rect 456 -107 462 -105
rect 450 -113 456 -111
rect 450 -115 452 -113
rect 454 -115 456 -113
rect 450 -117 456 -115
rect 450 -120 452 -117
rect 460 -120 462 -107
rect 470 -106 476 -104
rect 470 -108 472 -106
rect 474 -108 476 -106
rect 470 -110 476 -108
rect 480 -106 502 -104
rect 480 -108 491 -106
rect 493 -108 498 -106
rect 500 -108 502 -106
rect 480 -110 502 -108
rect 506 -106 512 -104
rect 506 -108 508 -106
rect 510 -108 512 -106
rect 506 -110 512 -108
rect 516 -106 522 -104
rect 516 -108 518 -106
rect 520 -108 522 -106
rect 516 -110 522 -108
rect 470 -113 472 -110
rect 480 -113 482 -110
rect 500 -113 502 -110
rect 507 -113 509 -110
rect 410 -128 412 -124
rect 420 -128 422 -124
rect 430 -128 432 -124
rect 371 -137 373 -133
rect 378 -137 380 -133
rect 389 -137 391 -133
rect 450 -137 452 -133
rect 460 -135 462 -130
rect 470 -132 472 -127
rect 480 -132 482 -127
rect 518 -119 520 -110
rect 539 -111 541 -98
rect 552 -101 554 -98
rect 641 -73 643 -69
rect 648 -73 650 -69
rect 628 -82 630 -78
rect 545 -103 554 -101
rect 545 -105 547 -103
rect 549 -105 551 -103
rect 562 -104 564 -101
rect 569 -104 571 -101
rect 587 -104 589 -101
rect 597 -104 599 -101
rect 607 -104 609 -101
rect 628 -103 630 -94
rect 641 -96 643 -91
rect 638 -98 644 -96
rect 638 -100 640 -98
rect 642 -100 644 -98
rect 638 -102 644 -100
rect 545 -107 551 -105
rect 539 -113 545 -111
rect 539 -115 541 -113
rect 543 -115 545 -113
rect 539 -117 545 -115
rect 539 -120 541 -117
rect 549 -120 551 -107
rect 559 -106 565 -104
rect 559 -108 561 -106
rect 563 -108 565 -106
rect 559 -110 565 -108
rect 569 -106 591 -104
rect 569 -108 580 -106
rect 582 -108 587 -106
rect 589 -108 591 -106
rect 569 -110 591 -108
rect 595 -106 601 -104
rect 595 -108 597 -106
rect 599 -108 601 -106
rect 595 -110 601 -108
rect 605 -106 611 -104
rect 605 -108 607 -106
rect 609 -108 611 -106
rect 605 -110 611 -108
rect 628 -105 634 -103
rect 628 -107 630 -105
rect 632 -107 634 -105
rect 628 -109 634 -107
rect 559 -113 561 -110
rect 569 -113 571 -110
rect 589 -113 591 -110
rect 596 -113 598 -110
rect 500 -137 502 -133
rect 507 -137 509 -133
rect 518 -137 520 -133
rect 539 -137 541 -133
rect 549 -135 551 -130
rect 559 -132 561 -127
rect 569 -132 571 -127
rect 607 -119 609 -110
rect 628 -118 630 -109
rect 638 -118 640 -102
rect 648 -104 650 -91
rect 648 -106 654 -104
rect 648 -108 650 -106
rect 652 -108 654 -106
rect 648 -110 654 -108
rect 648 -118 650 -110
rect 628 -128 630 -124
rect 638 -128 640 -124
rect 648 -128 650 -124
rect 589 -137 591 -133
rect 596 -137 598 -133
rect 607 -137 609 -133
rect 291 -145 293 -141
rect 302 -145 304 -141
rect 309 -145 311 -141
rect 239 -154 241 -150
rect 249 -154 251 -150
rect 259 -154 261 -150
rect 239 -168 241 -160
rect 235 -170 241 -168
rect 235 -172 237 -170
rect 239 -172 241 -170
rect 235 -174 241 -172
rect 239 -187 241 -174
rect 249 -176 251 -160
rect 259 -169 261 -160
rect 291 -168 293 -159
rect 329 -151 331 -146
rect 339 -151 341 -146
rect 349 -148 351 -143
rect 359 -145 361 -141
rect 391 -145 393 -141
rect 402 -145 404 -141
rect 409 -145 411 -141
rect 302 -168 304 -165
rect 309 -168 311 -165
rect 329 -168 331 -165
rect 339 -168 341 -165
rect 255 -171 261 -169
rect 255 -173 257 -171
rect 259 -173 261 -171
rect 255 -175 261 -173
rect 289 -170 295 -168
rect 289 -172 291 -170
rect 293 -172 295 -170
rect 289 -174 295 -172
rect 299 -170 305 -168
rect 299 -172 301 -170
rect 303 -172 305 -170
rect 299 -174 305 -172
rect 309 -170 331 -168
rect 309 -172 311 -170
rect 313 -172 318 -170
rect 320 -172 331 -170
rect 309 -174 331 -172
rect 335 -170 341 -168
rect 335 -172 337 -170
rect 339 -172 341 -170
rect 335 -174 341 -172
rect 349 -171 351 -158
rect 359 -161 361 -158
rect 355 -163 361 -161
rect 355 -165 357 -163
rect 359 -165 361 -163
rect 355 -167 361 -165
rect 349 -173 355 -171
rect 245 -178 251 -176
rect 245 -180 247 -178
rect 249 -180 251 -178
rect 245 -182 251 -180
rect 246 -187 248 -182
rect 259 -184 261 -175
rect 291 -177 293 -174
rect 301 -177 303 -174
rect 311 -177 313 -174
rect 329 -177 331 -174
rect 336 -177 338 -174
rect 349 -175 351 -173
rect 353 -175 355 -173
rect 346 -177 355 -175
rect 259 -200 261 -196
rect 239 -209 241 -205
rect 246 -209 248 -205
rect 346 -180 348 -177
rect 359 -180 361 -167
rect 391 -168 393 -159
rect 429 -151 431 -146
rect 439 -151 441 -146
rect 449 -148 451 -143
rect 459 -145 461 -141
rect 535 -145 537 -141
rect 546 -145 548 -141
rect 553 -145 555 -141
rect 483 -154 485 -150
rect 493 -154 495 -150
rect 503 -154 505 -150
rect 402 -168 404 -165
rect 409 -168 411 -165
rect 429 -168 431 -165
rect 439 -168 441 -165
rect 389 -170 395 -168
rect 389 -172 391 -170
rect 393 -172 395 -170
rect 389 -174 395 -172
rect 399 -170 405 -168
rect 399 -172 401 -170
rect 403 -172 405 -170
rect 399 -174 405 -172
rect 409 -170 431 -168
rect 409 -172 411 -170
rect 413 -172 418 -170
rect 420 -172 431 -170
rect 409 -174 431 -172
rect 435 -170 441 -168
rect 435 -172 437 -170
rect 439 -172 441 -170
rect 435 -174 441 -172
rect 449 -171 451 -158
rect 459 -161 461 -158
rect 455 -163 461 -161
rect 455 -165 457 -163
rect 459 -165 461 -163
rect 455 -167 461 -165
rect 449 -173 455 -171
rect 391 -177 393 -174
rect 401 -177 403 -174
rect 411 -177 413 -174
rect 429 -177 431 -174
rect 436 -177 438 -174
rect 449 -175 451 -173
rect 453 -175 455 -173
rect 446 -177 455 -175
rect 346 -198 348 -193
rect 291 -209 293 -205
rect 301 -209 303 -205
rect 311 -209 313 -205
rect 329 -207 331 -202
rect 336 -207 338 -202
rect 446 -180 448 -177
rect 459 -180 461 -167
rect 483 -168 485 -160
rect 479 -170 485 -168
rect 479 -172 481 -170
rect 483 -172 485 -170
rect 479 -174 485 -172
rect 446 -198 448 -193
rect 359 -209 361 -205
rect 391 -209 393 -205
rect 401 -209 403 -205
rect 411 -209 413 -205
rect 429 -207 431 -202
rect 436 -207 438 -202
rect 483 -187 485 -174
rect 493 -176 495 -160
rect 503 -169 505 -160
rect 535 -168 537 -159
rect 573 -151 575 -146
rect 583 -151 585 -146
rect 593 -148 595 -143
rect 603 -145 605 -141
rect 635 -145 637 -141
rect 646 -145 648 -141
rect 653 -145 655 -141
rect 546 -168 548 -165
rect 553 -168 555 -165
rect 573 -168 575 -165
rect 583 -168 585 -165
rect 499 -171 505 -169
rect 499 -173 501 -171
rect 503 -173 505 -171
rect 499 -175 505 -173
rect 533 -170 539 -168
rect 533 -172 535 -170
rect 537 -172 539 -170
rect 533 -174 539 -172
rect 543 -170 549 -168
rect 543 -172 545 -170
rect 547 -172 549 -170
rect 543 -174 549 -172
rect 553 -170 575 -168
rect 553 -172 555 -170
rect 557 -172 562 -170
rect 564 -172 575 -170
rect 553 -174 575 -172
rect 579 -170 585 -168
rect 579 -172 581 -170
rect 583 -172 585 -170
rect 579 -174 585 -172
rect 593 -171 595 -158
rect 603 -161 605 -158
rect 599 -163 605 -161
rect 599 -165 601 -163
rect 603 -165 605 -163
rect 599 -167 605 -165
rect 593 -173 599 -171
rect 489 -178 495 -176
rect 489 -180 491 -178
rect 493 -180 495 -178
rect 489 -182 495 -180
rect 490 -187 492 -182
rect 503 -184 505 -175
rect 535 -177 537 -174
rect 545 -177 547 -174
rect 555 -177 557 -174
rect 573 -177 575 -174
rect 580 -177 582 -174
rect 593 -175 595 -173
rect 597 -175 599 -173
rect 590 -177 599 -175
rect 503 -200 505 -196
rect 459 -209 461 -205
rect 483 -209 485 -205
rect 490 -209 492 -205
rect 590 -180 592 -177
rect 603 -180 605 -167
rect 635 -168 637 -159
rect 673 -151 675 -146
rect 683 -151 685 -146
rect 693 -148 695 -143
rect 703 -145 705 -141
rect 646 -168 648 -165
rect 653 -168 655 -165
rect 673 -168 675 -165
rect 683 -168 685 -165
rect 633 -170 639 -168
rect 633 -172 635 -170
rect 637 -172 639 -170
rect 633 -174 639 -172
rect 643 -170 649 -168
rect 643 -172 645 -170
rect 647 -172 649 -170
rect 643 -174 649 -172
rect 653 -170 675 -168
rect 653 -172 655 -170
rect 657 -172 662 -170
rect 664 -172 675 -170
rect 653 -174 675 -172
rect 679 -170 685 -168
rect 679 -172 681 -170
rect 683 -172 685 -170
rect 679 -174 685 -172
rect 693 -171 695 -158
rect 703 -161 705 -158
rect 699 -163 705 -161
rect 699 -165 701 -163
rect 703 -165 705 -163
rect 699 -167 705 -165
rect 693 -173 699 -171
rect 635 -177 637 -174
rect 645 -177 647 -174
rect 655 -177 657 -174
rect 673 -177 675 -174
rect 680 -177 682 -174
rect 693 -175 695 -173
rect 697 -175 699 -173
rect 690 -177 699 -175
rect 590 -198 592 -193
rect 535 -209 537 -205
rect 545 -209 547 -205
rect 555 -209 557 -205
rect 573 -207 575 -202
rect 580 -207 582 -202
rect 690 -180 692 -177
rect 703 -180 705 -167
rect 690 -198 692 -193
rect 603 -209 605 -205
rect 635 -209 637 -205
rect 645 -209 647 -205
rect 655 -209 657 -205
rect 673 -207 675 -202
rect 680 -207 682 -202
rect 703 -209 705 -205
rect 14 -217 16 -213
rect 37 -220 39 -215
rect 44 -220 46 -215
rect 62 -217 64 -213
rect 72 -217 74 -213
rect 82 -217 84 -213
rect 114 -217 116 -213
rect 27 -229 29 -224
rect 14 -255 16 -242
rect 27 -245 29 -242
rect 137 -220 139 -215
rect 144 -220 146 -215
rect 162 -217 164 -213
rect 172 -217 174 -213
rect 182 -217 184 -213
rect 127 -229 129 -224
rect 20 -247 29 -245
rect 20 -249 22 -247
rect 24 -249 26 -247
rect 37 -248 39 -245
rect 44 -248 46 -245
rect 62 -248 64 -245
rect 72 -248 74 -245
rect 82 -248 84 -245
rect 20 -251 26 -249
rect 14 -257 20 -255
rect 14 -259 16 -257
rect 18 -259 20 -257
rect 14 -261 20 -259
rect 14 -264 16 -261
rect 24 -264 26 -251
rect 34 -250 40 -248
rect 34 -252 36 -250
rect 38 -252 40 -250
rect 34 -254 40 -252
rect 44 -250 66 -248
rect 44 -252 55 -250
rect 57 -252 62 -250
rect 64 -252 66 -250
rect 44 -254 66 -252
rect 70 -250 76 -248
rect 70 -252 72 -250
rect 74 -252 76 -250
rect 70 -254 76 -252
rect 80 -250 86 -248
rect 80 -252 82 -250
rect 84 -252 86 -250
rect 80 -254 86 -252
rect 34 -257 36 -254
rect 44 -257 46 -254
rect 64 -257 66 -254
rect 71 -257 73 -254
rect 14 -281 16 -277
rect 24 -279 26 -274
rect 34 -276 36 -271
rect 44 -276 46 -271
rect 82 -263 84 -254
rect 114 -255 116 -242
rect 127 -245 129 -242
rect 227 -217 229 -213
rect 234 -217 236 -213
rect 255 -217 257 -213
rect 214 -226 216 -222
rect 120 -247 129 -245
rect 120 -249 122 -247
rect 124 -249 126 -247
rect 137 -248 139 -245
rect 144 -248 146 -245
rect 162 -248 164 -245
rect 172 -248 174 -245
rect 182 -248 184 -245
rect 214 -247 216 -238
rect 227 -240 229 -235
rect 224 -242 230 -240
rect 224 -244 226 -242
rect 228 -244 230 -242
rect 224 -246 230 -244
rect 120 -251 126 -249
rect 114 -257 120 -255
rect 114 -259 116 -257
rect 118 -259 120 -257
rect 114 -261 120 -259
rect 114 -264 116 -261
rect 124 -264 126 -251
rect 134 -250 140 -248
rect 134 -252 136 -250
rect 138 -252 140 -250
rect 134 -254 140 -252
rect 144 -250 166 -248
rect 144 -252 155 -250
rect 157 -252 162 -250
rect 164 -252 166 -250
rect 144 -254 166 -252
rect 170 -250 176 -248
rect 170 -252 172 -250
rect 174 -252 176 -250
rect 170 -254 176 -252
rect 180 -250 186 -248
rect 180 -252 182 -250
rect 184 -252 186 -250
rect 180 -254 186 -252
rect 214 -249 220 -247
rect 214 -251 216 -249
rect 218 -251 220 -249
rect 214 -253 220 -251
rect 134 -257 136 -254
rect 144 -257 146 -254
rect 164 -257 166 -254
rect 171 -257 173 -254
rect 64 -281 66 -277
rect 71 -281 73 -277
rect 82 -281 84 -277
rect 114 -281 116 -277
rect 124 -279 126 -274
rect 134 -276 136 -271
rect 144 -276 146 -271
rect 182 -263 184 -254
rect 214 -262 216 -253
rect 224 -262 226 -246
rect 234 -248 236 -235
rect 278 -220 280 -215
rect 285 -220 287 -215
rect 303 -217 305 -213
rect 313 -217 315 -213
rect 323 -217 325 -213
rect 355 -217 357 -213
rect 268 -229 270 -224
rect 234 -250 240 -248
rect 234 -252 236 -250
rect 238 -252 240 -250
rect 234 -254 240 -252
rect 234 -262 236 -254
rect 255 -255 257 -242
rect 268 -245 270 -242
rect 378 -220 380 -215
rect 385 -220 387 -215
rect 403 -217 405 -213
rect 413 -217 415 -213
rect 423 -217 425 -213
rect 368 -229 370 -224
rect 261 -247 270 -245
rect 261 -249 263 -247
rect 265 -249 267 -247
rect 278 -248 280 -245
rect 285 -248 287 -245
rect 303 -248 305 -245
rect 313 -248 315 -245
rect 323 -248 325 -245
rect 261 -251 267 -249
rect 255 -257 261 -255
rect 255 -259 257 -257
rect 259 -259 261 -257
rect 255 -261 261 -259
rect 255 -264 257 -261
rect 265 -264 267 -251
rect 275 -250 281 -248
rect 275 -252 277 -250
rect 279 -252 281 -250
rect 275 -254 281 -252
rect 285 -250 307 -248
rect 285 -252 296 -250
rect 298 -252 303 -250
rect 305 -252 307 -250
rect 285 -254 307 -252
rect 311 -250 317 -248
rect 311 -252 313 -250
rect 315 -252 317 -250
rect 311 -254 317 -252
rect 321 -250 327 -248
rect 321 -252 323 -250
rect 325 -252 327 -250
rect 321 -254 327 -252
rect 275 -257 277 -254
rect 285 -257 287 -254
rect 305 -257 307 -254
rect 312 -257 314 -254
rect 214 -272 216 -268
rect 224 -272 226 -268
rect 234 -272 236 -268
rect 164 -281 166 -277
rect 171 -281 173 -277
rect 182 -281 184 -277
rect 255 -281 257 -277
rect 265 -279 267 -274
rect 275 -276 277 -271
rect 285 -276 287 -271
rect 323 -263 325 -254
rect 355 -255 357 -242
rect 368 -245 370 -242
rect 468 -217 470 -213
rect 475 -217 477 -213
rect 455 -226 457 -222
rect 361 -247 370 -245
rect 361 -249 363 -247
rect 365 -249 367 -247
rect 378 -248 380 -245
rect 385 -248 387 -245
rect 403 -248 405 -245
rect 413 -248 415 -245
rect 423 -248 425 -245
rect 455 -247 457 -238
rect 468 -240 470 -235
rect 465 -242 471 -240
rect 465 -244 467 -242
rect 469 -244 471 -242
rect 465 -246 471 -244
rect 361 -251 367 -249
rect 355 -257 361 -255
rect 355 -259 357 -257
rect 359 -259 361 -257
rect 355 -261 361 -259
rect 355 -264 357 -261
rect 365 -264 367 -251
rect 375 -250 381 -248
rect 375 -252 377 -250
rect 379 -252 381 -250
rect 375 -254 381 -252
rect 385 -250 407 -248
rect 385 -252 396 -250
rect 398 -252 403 -250
rect 405 -252 407 -250
rect 385 -254 407 -252
rect 411 -250 417 -248
rect 411 -252 413 -250
rect 415 -252 417 -250
rect 411 -254 417 -252
rect 421 -250 427 -248
rect 421 -252 423 -250
rect 425 -252 427 -250
rect 421 -254 427 -252
rect 455 -249 461 -247
rect 455 -251 457 -249
rect 459 -251 461 -249
rect 455 -253 461 -251
rect 375 -257 377 -254
rect 385 -257 387 -254
rect 405 -257 407 -254
rect 412 -257 414 -254
rect 305 -281 307 -277
rect 312 -281 314 -277
rect 323 -281 325 -277
rect 355 -281 357 -277
rect 365 -279 367 -274
rect 375 -276 377 -271
rect 385 -276 387 -271
rect 423 -263 425 -254
rect 455 -262 457 -253
rect 465 -262 467 -246
rect 475 -248 477 -235
rect 475 -250 481 -248
rect 475 -252 477 -250
rect 479 -252 481 -250
rect 475 -254 481 -252
rect 475 -262 477 -254
rect 455 -272 457 -268
rect 465 -272 467 -268
rect 475 -272 477 -268
rect 405 -281 407 -277
rect 412 -281 414 -277
rect 423 -281 425 -277
<< ndif >>
rect 7 24 14 26
rect 7 22 9 24
rect 11 22 14 24
rect 7 20 14 22
rect 16 23 24 26
rect 51 24 58 26
rect 16 20 26 23
rect 18 14 26 20
rect 28 14 33 23
rect 35 21 42 23
rect 35 19 38 21
rect 40 19 42 21
rect 51 22 53 24
rect 55 22 58 24
rect 51 20 58 22
rect 60 23 68 26
rect 95 24 102 26
rect 60 20 70 23
rect 35 17 42 19
rect 35 14 40 17
rect 62 14 70 20
rect 72 14 77 23
rect 79 21 86 23
rect 79 19 82 21
rect 84 19 86 21
rect 95 22 97 24
rect 99 22 102 24
rect 95 20 102 22
rect 104 23 112 26
rect 139 24 146 26
rect 104 20 114 23
rect 79 17 86 19
rect 79 14 84 17
rect 106 14 114 20
rect 116 14 121 23
rect 123 21 130 23
rect 123 19 126 21
rect 128 19 130 21
rect 139 22 141 24
rect 143 22 146 24
rect 139 20 146 22
rect 148 23 156 26
rect 183 24 190 26
rect 148 20 158 23
rect 123 17 130 19
rect 123 14 128 17
rect 150 14 158 20
rect 160 14 165 23
rect 167 21 174 23
rect 167 19 170 21
rect 172 19 174 21
rect 183 22 185 24
rect 187 22 190 24
rect 183 20 190 22
rect 192 23 200 26
rect 227 24 234 26
rect 192 20 202 23
rect 167 17 174 19
rect 167 14 172 17
rect 194 14 202 20
rect 204 14 209 23
rect 211 21 218 23
rect 211 19 214 21
rect 216 19 218 21
rect 227 22 229 24
rect 231 22 234 24
rect 227 20 234 22
rect 236 23 244 26
rect 271 24 278 26
rect 236 20 246 23
rect 211 17 218 19
rect 211 14 216 17
rect 238 14 246 20
rect 248 14 253 23
rect 255 21 262 23
rect 255 19 258 21
rect 260 19 262 21
rect 271 22 273 24
rect 275 22 278 24
rect 271 20 278 22
rect 280 23 288 26
rect 315 24 322 26
rect 280 20 290 23
rect 255 17 262 19
rect 255 14 260 17
rect 282 14 290 20
rect 292 14 297 23
rect 299 21 306 23
rect 299 19 302 21
rect 304 19 306 21
rect 315 22 317 24
rect 319 22 322 24
rect 315 20 322 22
rect 324 23 332 26
rect 359 24 366 26
rect 324 20 334 23
rect 299 17 306 19
rect 299 14 304 17
rect 326 14 334 20
rect 336 14 341 23
rect 343 21 350 23
rect 343 19 346 21
rect 348 19 350 21
rect 359 22 361 24
rect 363 22 366 24
rect 359 20 366 22
rect 368 23 376 26
rect 403 24 410 26
rect 368 20 378 23
rect 343 17 350 19
rect 343 14 348 17
rect 370 14 378 20
rect 380 14 385 23
rect 387 21 394 23
rect 387 19 390 21
rect 392 19 394 21
rect 403 22 405 24
rect 407 22 410 24
rect 403 20 410 22
rect 412 23 420 26
rect 447 24 454 26
rect 412 20 422 23
rect 387 17 394 19
rect 387 14 392 17
rect 414 14 422 20
rect 424 14 429 23
rect 431 21 438 23
rect 431 19 434 21
rect 436 19 438 21
rect 447 22 449 24
rect 451 22 454 24
rect 447 20 454 22
rect 456 23 464 26
rect 491 24 498 26
rect 456 20 466 23
rect 431 17 438 19
rect 431 14 436 17
rect 458 14 466 20
rect 468 14 473 23
rect 475 21 482 23
rect 475 19 478 21
rect 480 19 482 21
rect 491 22 493 24
rect 495 22 498 24
rect 491 20 498 22
rect 500 23 508 26
rect 535 24 542 26
rect 500 20 510 23
rect 475 17 482 19
rect 475 14 480 17
rect 502 14 510 20
rect 512 14 517 23
rect 519 21 526 23
rect 519 19 522 21
rect 524 19 526 21
rect 535 22 537 24
rect 539 22 542 24
rect 535 20 542 22
rect 544 23 552 26
rect 579 24 586 26
rect 544 20 554 23
rect 519 17 526 19
rect 519 14 524 17
rect 546 14 554 20
rect 556 14 561 23
rect 563 21 570 23
rect 563 19 566 21
rect 568 19 570 21
rect 579 22 581 24
rect 583 22 586 24
rect 579 20 586 22
rect 588 23 596 26
rect 623 24 630 26
rect 588 20 598 23
rect 563 17 570 19
rect 563 14 568 17
rect 590 14 598 20
rect 600 14 605 23
rect 607 21 614 23
rect 607 19 610 21
rect 612 19 614 21
rect 623 22 625 24
rect 627 22 630 24
rect 623 20 630 22
rect 632 23 640 26
rect 667 24 674 26
rect 632 20 642 23
rect 607 17 614 19
rect 607 14 612 17
rect 634 14 642 20
rect 644 14 649 23
rect 651 21 658 23
rect 651 19 654 21
rect 656 19 658 21
rect 667 22 669 24
rect 671 22 674 24
rect 667 20 674 22
rect 676 23 684 26
rect 676 20 686 23
rect 651 17 658 19
rect 651 14 656 17
rect 678 14 686 20
rect 688 14 693 23
rect 695 21 702 23
rect 695 19 698 21
rect 700 19 702 21
rect 695 17 702 19
rect 695 14 700 17
rect 18 12 24 14
rect 18 10 20 12
rect 22 10 24 12
rect 18 8 24 10
rect 62 12 68 14
rect 62 10 64 12
rect 66 10 68 12
rect 62 8 68 10
rect 106 12 112 14
rect 106 10 108 12
rect 110 10 112 12
rect 106 8 112 10
rect 150 12 156 14
rect 150 10 152 12
rect 154 10 156 12
rect 150 8 156 10
rect 194 12 200 14
rect 194 10 196 12
rect 198 10 200 12
rect 194 8 200 10
rect 238 12 244 14
rect 238 10 240 12
rect 242 10 244 12
rect 238 8 244 10
rect 282 12 288 14
rect 282 10 284 12
rect 286 10 288 12
rect 282 8 288 10
rect 326 12 332 14
rect 326 10 328 12
rect 330 10 332 12
rect 326 8 332 10
rect 370 12 376 14
rect 370 10 372 12
rect 374 10 376 12
rect 370 8 376 10
rect 414 12 420 14
rect 414 10 416 12
rect 418 10 420 12
rect 414 8 420 10
rect 458 12 464 14
rect 458 10 460 12
rect 462 10 464 12
rect 458 8 464 10
rect 502 12 508 14
rect 502 10 504 12
rect 506 10 508 12
rect 502 8 508 10
rect 546 12 552 14
rect 546 10 548 12
rect 550 10 552 12
rect 546 8 552 10
rect 590 12 596 14
rect 590 10 592 12
rect 594 10 596 12
rect 590 8 596 10
rect 634 12 640 14
rect 634 10 636 12
rect 638 10 640 12
rect 634 8 640 10
rect 678 12 684 14
rect 678 10 680 12
rect 682 10 684 12
rect 678 8 684 10
rect 17 -8 22 -1
rect 15 -10 22 -8
rect 15 -12 17 -10
rect 19 -12 22 -10
rect 15 -15 22 -12
rect 24 -3 33 -1
rect 24 -5 28 -3
rect 30 -5 33 -3
rect 24 -15 33 -5
rect 26 -21 33 -15
rect 35 -21 40 -1
rect 42 -8 47 -1
rect 85 -4 90 -1
rect 75 -7 80 -4
rect 42 -10 49 -8
rect 42 -12 45 -10
rect 47 -12 49 -10
rect 42 -14 49 -12
rect 53 -10 60 -7
rect 53 -12 55 -10
rect 57 -12 60 -10
rect 42 -21 47 -14
rect 53 -17 60 -12
rect 53 -19 55 -17
rect 57 -19 60 -17
rect 53 -21 60 -19
rect 62 -17 70 -7
rect 62 -19 65 -17
rect 67 -19 70 -17
rect 62 -21 70 -19
rect 72 -9 80 -7
rect 72 -11 75 -9
rect 77 -11 80 -9
rect 72 -14 80 -11
rect 82 -6 90 -4
rect 82 -8 85 -6
rect 87 -8 90 -6
rect 82 -14 90 -8
rect 92 -8 97 -1
rect 106 -8 111 -1
rect 92 -10 99 -8
rect 92 -12 95 -10
rect 97 -12 99 -10
rect 92 -14 99 -12
rect 104 -10 111 -8
rect 104 -12 106 -10
rect 108 -12 111 -10
rect 72 -21 77 -14
rect 104 -15 111 -12
rect 113 -3 122 -1
rect 113 -5 117 -3
rect 119 -5 122 -3
rect 113 -15 122 -5
rect 115 -21 122 -15
rect 124 -21 129 -1
rect 131 -8 136 -1
rect 174 -4 179 -1
rect 164 -7 169 -4
rect 131 -10 138 -8
rect 131 -12 134 -10
rect 136 -12 138 -10
rect 131 -14 138 -12
rect 142 -10 149 -7
rect 142 -12 144 -10
rect 146 -12 149 -10
rect 131 -21 136 -14
rect 142 -17 149 -12
rect 142 -19 144 -17
rect 146 -19 149 -17
rect 142 -21 149 -19
rect 151 -17 159 -7
rect 151 -19 154 -17
rect 156 -19 159 -17
rect 151 -21 159 -19
rect 161 -9 169 -7
rect 161 -11 164 -9
rect 166 -11 169 -9
rect 161 -14 169 -11
rect 171 -6 179 -4
rect 171 -8 174 -6
rect 176 -8 179 -6
rect 171 -14 179 -8
rect 181 -8 186 -1
rect 181 -10 188 -8
rect 235 -8 240 -1
rect 233 -10 240 -8
rect 181 -12 184 -10
rect 186 -12 188 -10
rect 181 -14 188 -12
rect 192 -12 199 -10
rect 192 -14 194 -12
rect 196 -14 199 -12
rect 161 -21 166 -14
rect 192 -16 199 -14
rect 201 -12 209 -10
rect 201 -14 204 -12
rect 206 -14 209 -12
rect 201 -16 209 -14
rect 211 -12 219 -10
rect 211 -14 214 -12
rect 216 -14 219 -12
rect 211 -16 219 -14
rect 221 -12 228 -10
rect 221 -14 224 -12
rect 226 -14 228 -12
rect 221 -16 228 -14
rect 233 -12 235 -10
rect 237 -12 240 -10
rect 233 -15 240 -12
rect 242 -3 251 -1
rect 242 -5 246 -3
rect 248 -5 251 -3
rect 242 -15 251 -5
rect 244 -21 251 -15
rect 253 -21 258 -1
rect 260 -8 265 -1
rect 303 -4 308 -1
rect 293 -7 298 -4
rect 260 -10 267 -8
rect 260 -12 263 -10
rect 265 -12 267 -10
rect 260 -14 267 -12
rect 271 -10 278 -7
rect 271 -12 273 -10
rect 275 -12 278 -10
rect 260 -21 265 -14
rect 271 -17 278 -12
rect 271 -19 273 -17
rect 275 -19 278 -17
rect 271 -21 278 -19
rect 280 -17 288 -7
rect 280 -19 283 -17
rect 285 -19 288 -17
rect 280 -21 288 -19
rect 290 -9 298 -7
rect 290 -11 293 -9
rect 295 -11 298 -9
rect 290 -14 298 -11
rect 300 -6 308 -4
rect 300 -8 303 -6
rect 305 -8 308 -6
rect 300 -14 308 -8
rect 310 -8 315 -1
rect 324 -8 329 -1
rect 310 -10 317 -8
rect 310 -12 313 -10
rect 315 -12 317 -10
rect 310 -14 317 -12
rect 322 -10 329 -8
rect 322 -12 324 -10
rect 326 -12 329 -10
rect 290 -21 295 -14
rect 322 -15 329 -12
rect 331 -3 340 -1
rect 331 -5 335 -3
rect 337 -5 340 -3
rect 331 -15 340 -5
rect 333 -21 340 -15
rect 342 -21 347 -1
rect 349 -8 354 -1
rect 392 -4 397 -1
rect 382 -7 387 -4
rect 349 -10 356 -8
rect 349 -12 352 -10
rect 354 -12 356 -10
rect 349 -14 356 -12
rect 360 -10 367 -7
rect 360 -12 362 -10
rect 364 -12 367 -10
rect 349 -21 354 -14
rect 360 -17 367 -12
rect 360 -19 362 -17
rect 364 -19 367 -17
rect 360 -21 367 -19
rect 369 -17 377 -7
rect 369 -19 372 -17
rect 374 -19 377 -17
rect 369 -21 377 -19
rect 379 -9 387 -7
rect 379 -11 382 -9
rect 384 -11 387 -9
rect 379 -14 387 -11
rect 389 -6 397 -4
rect 389 -8 392 -6
rect 394 -8 397 -6
rect 389 -14 397 -8
rect 399 -8 404 -1
rect 493 -8 498 -1
rect 399 -10 406 -8
rect 399 -12 402 -10
rect 404 -12 406 -10
rect 399 -14 406 -12
rect 491 -10 498 -8
rect 491 -12 493 -10
rect 495 -12 498 -10
rect 379 -21 384 -14
rect 491 -15 498 -12
rect 500 -3 509 -1
rect 500 -5 504 -3
rect 506 -5 509 -3
rect 500 -15 509 -5
rect 502 -21 509 -15
rect 511 -21 516 -1
rect 518 -8 523 -1
rect 561 -4 566 -1
rect 551 -7 556 -4
rect 518 -10 525 -8
rect 518 -12 521 -10
rect 523 -12 525 -10
rect 518 -14 525 -12
rect 529 -10 536 -7
rect 529 -12 531 -10
rect 533 -12 536 -10
rect 518 -21 523 -14
rect 529 -17 536 -12
rect 529 -19 531 -17
rect 533 -19 536 -17
rect 529 -21 536 -19
rect 538 -17 546 -7
rect 538 -19 541 -17
rect 543 -19 546 -17
rect 538 -21 546 -19
rect 548 -9 556 -7
rect 548 -11 551 -9
rect 553 -11 556 -9
rect 548 -14 556 -11
rect 558 -6 566 -4
rect 558 -8 561 -6
rect 563 -8 566 -6
rect 558 -14 566 -8
rect 568 -8 573 -1
rect 582 -8 587 -1
rect 568 -10 575 -8
rect 568 -12 571 -10
rect 573 -12 575 -10
rect 568 -14 575 -12
rect 580 -10 587 -8
rect 580 -12 582 -10
rect 584 -12 587 -10
rect 548 -21 553 -14
rect 580 -15 587 -12
rect 589 -3 598 -1
rect 589 -5 593 -3
rect 595 -5 598 -3
rect 589 -15 598 -5
rect 591 -21 598 -15
rect 600 -21 605 -1
rect 607 -8 612 -1
rect 650 -4 655 -1
rect 640 -7 645 -4
rect 607 -10 614 -8
rect 607 -12 610 -10
rect 612 -12 614 -10
rect 607 -14 614 -12
rect 618 -10 625 -7
rect 618 -12 620 -10
rect 622 -12 625 -10
rect 607 -21 612 -14
rect 618 -17 625 -12
rect 618 -19 620 -17
rect 622 -19 625 -17
rect 618 -21 625 -19
rect 627 -17 635 -7
rect 627 -19 630 -17
rect 632 -19 635 -17
rect 627 -21 635 -19
rect 637 -9 645 -7
rect 637 -11 640 -9
rect 642 -11 645 -9
rect 637 -14 645 -11
rect 647 -6 655 -4
rect 647 -8 650 -6
rect 652 -8 655 -6
rect 647 -14 655 -8
rect 657 -8 662 -1
rect 657 -10 664 -8
rect 657 -12 660 -10
rect 662 -12 664 -10
rect 657 -14 664 -12
rect 637 -21 642 -14
rect 29 -120 34 -113
rect 7 -122 14 -120
rect 7 -124 9 -122
rect 11 -124 14 -122
rect 7 -126 14 -124
rect 9 -133 14 -126
rect 16 -126 24 -120
rect 16 -128 19 -126
rect 21 -128 24 -126
rect 16 -130 24 -128
rect 26 -123 34 -120
rect 26 -125 29 -123
rect 31 -125 34 -123
rect 26 -127 34 -125
rect 36 -115 44 -113
rect 36 -117 39 -115
rect 41 -117 44 -115
rect 36 -127 44 -117
rect 46 -115 53 -113
rect 46 -117 49 -115
rect 51 -117 53 -115
rect 46 -122 53 -117
rect 59 -120 64 -113
rect 46 -124 49 -122
rect 51 -124 53 -122
rect 46 -127 53 -124
rect 57 -122 64 -120
rect 57 -124 59 -122
rect 61 -124 64 -122
rect 57 -126 64 -124
rect 26 -130 31 -127
rect 16 -133 21 -130
rect 59 -133 64 -126
rect 66 -133 71 -113
rect 73 -119 80 -113
rect 73 -129 82 -119
rect 73 -131 76 -129
rect 78 -131 82 -129
rect 73 -133 82 -131
rect 84 -122 91 -119
rect 118 -120 123 -113
rect 84 -124 87 -122
rect 89 -124 91 -122
rect 84 -126 91 -124
rect 96 -122 103 -120
rect 96 -124 98 -122
rect 100 -124 103 -122
rect 96 -126 103 -124
rect 84 -133 89 -126
rect 98 -133 103 -126
rect 105 -126 113 -120
rect 105 -128 108 -126
rect 110 -128 113 -126
rect 105 -130 113 -128
rect 115 -123 123 -120
rect 115 -125 118 -123
rect 120 -125 123 -123
rect 115 -127 123 -125
rect 125 -115 133 -113
rect 125 -117 128 -115
rect 130 -117 133 -115
rect 125 -127 133 -117
rect 135 -115 142 -113
rect 135 -117 138 -115
rect 140 -117 142 -115
rect 135 -122 142 -117
rect 148 -120 153 -113
rect 135 -124 138 -122
rect 140 -124 142 -122
rect 135 -127 142 -124
rect 146 -122 153 -120
rect 146 -124 148 -122
rect 150 -124 153 -122
rect 146 -126 153 -124
rect 115 -130 120 -127
rect 105 -133 110 -130
rect 148 -133 153 -126
rect 155 -133 160 -113
rect 162 -119 169 -113
rect 162 -129 171 -119
rect 162 -131 165 -129
rect 167 -131 171 -129
rect 162 -133 171 -131
rect 173 -122 180 -119
rect 173 -124 176 -122
rect 178 -124 180 -122
rect 185 -120 192 -118
rect 185 -122 187 -120
rect 189 -122 192 -120
rect 185 -124 192 -122
rect 194 -120 202 -118
rect 194 -122 197 -120
rect 199 -122 202 -120
rect 194 -124 202 -122
rect 204 -120 212 -118
rect 204 -122 207 -120
rect 209 -122 212 -120
rect 204 -124 212 -122
rect 214 -120 221 -118
rect 247 -120 252 -113
rect 214 -122 217 -120
rect 219 -122 221 -120
rect 214 -124 221 -122
rect 225 -122 232 -120
rect 225 -124 227 -122
rect 229 -124 232 -122
rect 173 -126 180 -124
rect 173 -133 178 -126
rect 225 -126 232 -124
rect 227 -133 232 -126
rect 234 -126 242 -120
rect 234 -128 237 -126
rect 239 -128 242 -126
rect 234 -130 242 -128
rect 244 -123 252 -120
rect 244 -125 247 -123
rect 249 -125 252 -123
rect 244 -127 252 -125
rect 254 -115 262 -113
rect 254 -117 257 -115
rect 259 -117 262 -115
rect 254 -127 262 -117
rect 264 -115 271 -113
rect 264 -117 267 -115
rect 269 -117 271 -115
rect 264 -122 271 -117
rect 277 -120 282 -113
rect 264 -124 267 -122
rect 269 -124 271 -122
rect 264 -127 271 -124
rect 275 -122 282 -120
rect 275 -124 277 -122
rect 279 -124 282 -122
rect 275 -126 282 -124
rect 244 -130 249 -127
rect 234 -133 239 -130
rect 277 -133 282 -126
rect 284 -133 289 -113
rect 291 -119 298 -113
rect 291 -129 300 -119
rect 291 -131 294 -129
rect 296 -131 300 -129
rect 291 -133 300 -131
rect 302 -122 309 -119
rect 336 -120 341 -113
rect 302 -124 305 -122
rect 307 -124 309 -122
rect 302 -126 309 -124
rect 314 -122 321 -120
rect 314 -124 316 -122
rect 318 -124 321 -122
rect 314 -126 321 -124
rect 302 -133 307 -126
rect 316 -133 321 -126
rect 323 -126 331 -120
rect 323 -128 326 -126
rect 328 -128 331 -126
rect 323 -130 331 -128
rect 333 -123 341 -120
rect 333 -125 336 -123
rect 338 -125 341 -123
rect 333 -127 341 -125
rect 343 -115 351 -113
rect 343 -117 346 -115
rect 348 -117 351 -115
rect 343 -127 351 -117
rect 353 -115 360 -113
rect 353 -117 356 -115
rect 358 -117 360 -115
rect 353 -122 360 -117
rect 366 -120 371 -113
rect 353 -124 356 -122
rect 358 -124 360 -122
rect 353 -127 360 -124
rect 364 -122 371 -120
rect 364 -124 366 -122
rect 368 -124 371 -122
rect 364 -126 371 -124
rect 333 -130 338 -127
rect 323 -133 328 -130
rect 366 -133 371 -126
rect 373 -133 378 -113
rect 380 -119 387 -113
rect 380 -129 389 -119
rect 380 -131 383 -129
rect 385 -131 389 -129
rect 380 -133 389 -131
rect 391 -122 398 -119
rect 391 -124 394 -122
rect 396 -124 398 -122
rect 403 -120 410 -118
rect 403 -122 405 -120
rect 407 -122 410 -120
rect 403 -124 410 -122
rect 412 -120 420 -118
rect 412 -122 415 -120
rect 417 -122 420 -120
rect 412 -124 420 -122
rect 422 -120 430 -118
rect 422 -122 425 -120
rect 427 -122 430 -120
rect 422 -124 430 -122
rect 432 -120 439 -118
rect 465 -120 470 -113
rect 432 -122 435 -120
rect 437 -122 439 -120
rect 432 -124 439 -122
rect 443 -122 450 -120
rect 443 -124 445 -122
rect 447 -124 450 -122
rect 391 -126 398 -124
rect 391 -133 396 -126
rect 443 -126 450 -124
rect 445 -133 450 -126
rect 452 -126 460 -120
rect 452 -128 455 -126
rect 457 -128 460 -126
rect 452 -130 460 -128
rect 462 -123 470 -120
rect 462 -125 465 -123
rect 467 -125 470 -123
rect 462 -127 470 -125
rect 472 -115 480 -113
rect 472 -117 475 -115
rect 477 -117 480 -115
rect 472 -127 480 -117
rect 482 -115 489 -113
rect 482 -117 485 -115
rect 487 -117 489 -115
rect 482 -122 489 -117
rect 495 -120 500 -113
rect 482 -124 485 -122
rect 487 -124 489 -122
rect 482 -127 489 -124
rect 493 -122 500 -120
rect 493 -124 495 -122
rect 497 -124 500 -122
rect 493 -126 500 -124
rect 462 -130 467 -127
rect 452 -133 457 -130
rect 495 -133 500 -126
rect 502 -133 507 -113
rect 509 -119 516 -113
rect 509 -129 518 -119
rect 509 -131 512 -129
rect 514 -131 518 -129
rect 509 -133 518 -131
rect 520 -122 527 -119
rect 554 -120 559 -113
rect 520 -124 523 -122
rect 525 -124 527 -122
rect 520 -126 527 -124
rect 532 -122 539 -120
rect 532 -124 534 -122
rect 536 -124 539 -122
rect 532 -126 539 -124
rect 520 -133 525 -126
rect 534 -133 539 -126
rect 541 -126 549 -120
rect 541 -128 544 -126
rect 546 -128 549 -126
rect 541 -130 549 -128
rect 551 -123 559 -120
rect 551 -125 554 -123
rect 556 -125 559 -123
rect 551 -127 559 -125
rect 561 -115 569 -113
rect 561 -117 564 -115
rect 566 -117 569 -115
rect 561 -127 569 -117
rect 571 -115 578 -113
rect 571 -117 574 -115
rect 576 -117 578 -115
rect 571 -122 578 -117
rect 584 -120 589 -113
rect 571 -124 574 -122
rect 576 -124 578 -122
rect 571 -127 578 -124
rect 582 -122 589 -120
rect 582 -124 584 -122
rect 586 -124 589 -122
rect 582 -126 589 -124
rect 551 -130 556 -127
rect 541 -133 546 -130
rect 584 -133 589 -126
rect 591 -133 596 -113
rect 598 -119 605 -113
rect 598 -129 607 -119
rect 598 -131 601 -129
rect 603 -131 607 -129
rect 598 -133 607 -131
rect 609 -122 616 -119
rect 609 -124 612 -122
rect 614 -124 616 -122
rect 621 -120 628 -118
rect 621 -122 623 -120
rect 625 -122 628 -120
rect 621 -124 628 -122
rect 630 -120 638 -118
rect 630 -122 633 -120
rect 635 -122 638 -120
rect 630 -124 638 -122
rect 640 -120 648 -118
rect 640 -122 643 -120
rect 645 -122 648 -120
rect 640 -124 648 -122
rect 650 -120 657 -118
rect 650 -122 653 -120
rect 655 -122 657 -120
rect 650 -124 657 -122
rect 609 -126 616 -124
rect 609 -133 614 -126
rect 286 -152 291 -145
rect 284 -154 291 -152
rect 232 -156 239 -154
rect 232 -158 234 -156
rect 236 -158 239 -156
rect 232 -160 239 -158
rect 241 -156 249 -154
rect 241 -158 244 -156
rect 246 -158 249 -156
rect 241 -160 249 -158
rect 251 -156 259 -154
rect 251 -158 254 -156
rect 256 -158 259 -156
rect 251 -160 259 -158
rect 261 -156 268 -154
rect 261 -158 264 -156
rect 266 -158 268 -156
rect 261 -160 268 -158
rect 284 -156 286 -154
rect 288 -156 291 -154
rect 284 -159 291 -156
rect 293 -147 302 -145
rect 293 -149 297 -147
rect 299 -149 302 -147
rect 293 -159 302 -149
rect 295 -165 302 -159
rect 304 -165 309 -145
rect 311 -152 316 -145
rect 354 -148 359 -145
rect 344 -151 349 -148
rect 311 -154 318 -152
rect 311 -156 314 -154
rect 316 -156 318 -154
rect 311 -158 318 -156
rect 322 -154 329 -151
rect 322 -156 324 -154
rect 326 -156 329 -154
rect 311 -165 316 -158
rect 322 -161 329 -156
rect 322 -163 324 -161
rect 326 -163 329 -161
rect 322 -165 329 -163
rect 331 -161 339 -151
rect 331 -163 334 -161
rect 336 -163 339 -161
rect 331 -165 339 -163
rect 341 -153 349 -151
rect 341 -155 344 -153
rect 346 -155 349 -153
rect 341 -158 349 -155
rect 351 -150 359 -148
rect 351 -152 354 -150
rect 356 -152 359 -150
rect 351 -158 359 -152
rect 361 -152 366 -145
rect 386 -152 391 -145
rect 361 -154 368 -152
rect 361 -156 364 -154
rect 366 -156 368 -154
rect 361 -158 368 -156
rect 384 -154 391 -152
rect 384 -156 386 -154
rect 388 -156 391 -154
rect 341 -165 346 -158
rect 384 -159 391 -156
rect 393 -147 402 -145
rect 393 -149 397 -147
rect 399 -149 402 -147
rect 393 -159 402 -149
rect 395 -165 402 -159
rect 404 -165 409 -145
rect 411 -152 416 -145
rect 454 -148 459 -145
rect 444 -151 449 -148
rect 411 -154 418 -152
rect 411 -156 414 -154
rect 416 -156 418 -154
rect 411 -158 418 -156
rect 422 -154 429 -151
rect 422 -156 424 -154
rect 426 -156 429 -154
rect 411 -165 416 -158
rect 422 -161 429 -156
rect 422 -163 424 -161
rect 426 -163 429 -161
rect 422 -165 429 -163
rect 431 -161 439 -151
rect 431 -163 434 -161
rect 436 -163 439 -161
rect 431 -165 439 -163
rect 441 -153 449 -151
rect 441 -155 444 -153
rect 446 -155 449 -153
rect 441 -158 449 -155
rect 451 -150 459 -148
rect 451 -152 454 -150
rect 456 -152 459 -150
rect 451 -158 459 -152
rect 461 -152 466 -145
rect 461 -154 468 -152
rect 530 -152 535 -145
rect 528 -154 535 -152
rect 461 -156 464 -154
rect 466 -156 468 -154
rect 461 -158 468 -156
rect 476 -156 483 -154
rect 476 -158 478 -156
rect 480 -158 483 -156
rect 441 -165 446 -158
rect 476 -160 483 -158
rect 485 -156 493 -154
rect 485 -158 488 -156
rect 490 -158 493 -156
rect 485 -160 493 -158
rect 495 -156 503 -154
rect 495 -158 498 -156
rect 500 -158 503 -156
rect 495 -160 503 -158
rect 505 -156 512 -154
rect 505 -158 508 -156
rect 510 -158 512 -156
rect 505 -160 512 -158
rect 528 -156 530 -154
rect 532 -156 535 -154
rect 528 -159 535 -156
rect 537 -147 546 -145
rect 537 -149 541 -147
rect 543 -149 546 -147
rect 537 -159 546 -149
rect 539 -165 546 -159
rect 548 -165 553 -145
rect 555 -152 560 -145
rect 598 -148 603 -145
rect 588 -151 593 -148
rect 555 -154 562 -152
rect 555 -156 558 -154
rect 560 -156 562 -154
rect 555 -158 562 -156
rect 566 -154 573 -151
rect 566 -156 568 -154
rect 570 -156 573 -154
rect 555 -165 560 -158
rect 566 -161 573 -156
rect 566 -163 568 -161
rect 570 -163 573 -161
rect 566 -165 573 -163
rect 575 -161 583 -151
rect 575 -163 578 -161
rect 580 -163 583 -161
rect 575 -165 583 -163
rect 585 -153 593 -151
rect 585 -155 588 -153
rect 590 -155 593 -153
rect 585 -158 593 -155
rect 595 -150 603 -148
rect 595 -152 598 -150
rect 600 -152 603 -150
rect 595 -158 603 -152
rect 605 -152 610 -145
rect 630 -152 635 -145
rect 605 -154 612 -152
rect 605 -156 608 -154
rect 610 -156 612 -154
rect 605 -158 612 -156
rect 628 -154 635 -152
rect 628 -156 630 -154
rect 632 -156 635 -154
rect 585 -165 590 -158
rect 628 -159 635 -156
rect 637 -147 646 -145
rect 637 -149 641 -147
rect 643 -149 646 -147
rect 637 -159 646 -149
rect 639 -165 646 -159
rect 648 -165 653 -145
rect 655 -152 660 -145
rect 698 -148 703 -145
rect 688 -151 693 -148
rect 655 -154 662 -152
rect 655 -156 658 -154
rect 660 -156 662 -154
rect 655 -158 662 -156
rect 666 -154 673 -151
rect 666 -156 668 -154
rect 670 -156 673 -154
rect 655 -165 660 -158
rect 666 -161 673 -156
rect 666 -163 668 -161
rect 670 -163 673 -161
rect 666 -165 673 -163
rect 675 -161 683 -151
rect 675 -163 678 -161
rect 680 -163 683 -161
rect 675 -165 683 -163
rect 685 -153 693 -151
rect 685 -155 688 -153
rect 690 -155 693 -153
rect 685 -158 693 -155
rect 695 -150 703 -148
rect 695 -152 698 -150
rect 700 -152 703 -150
rect 695 -158 703 -152
rect 705 -152 710 -145
rect 705 -154 712 -152
rect 705 -156 708 -154
rect 710 -156 712 -154
rect 705 -158 712 -156
rect 685 -165 690 -158
rect 29 -264 34 -257
rect 7 -266 14 -264
rect 7 -268 9 -266
rect 11 -268 14 -266
rect 7 -270 14 -268
rect 9 -277 14 -270
rect 16 -270 24 -264
rect 16 -272 19 -270
rect 21 -272 24 -270
rect 16 -274 24 -272
rect 26 -267 34 -264
rect 26 -269 29 -267
rect 31 -269 34 -267
rect 26 -271 34 -269
rect 36 -259 44 -257
rect 36 -261 39 -259
rect 41 -261 44 -259
rect 36 -271 44 -261
rect 46 -259 53 -257
rect 46 -261 49 -259
rect 51 -261 53 -259
rect 46 -266 53 -261
rect 59 -264 64 -257
rect 46 -268 49 -266
rect 51 -268 53 -266
rect 46 -271 53 -268
rect 57 -266 64 -264
rect 57 -268 59 -266
rect 61 -268 64 -266
rect 57 -270 64 -268
rect 26 -274 31 -271
rect 16 -277 21 -274
rect 59 -277 64 -270
rect 66 -277 71 -257
rect 73 -263 80 -257
rect 73 -273 82 -263
rect 73 -275 76 -273
rect 78 -275 82 -273
rect 73 -277 82 -275
rect 84 -266 91 -263
rect 129 -264 134 -257
rect 84 -268 87 -266
rect 89 -268 91 -266
rect 84 -270 91 -268
rect 107 -266 114 -264
rect 107 -268 109 -266
rect 111 -268 114 -266
rect 107 -270 114 -268
rect 84 -277 89 -270
rect 109 -277 114 -270
rect 116 -270 124 -264
rect 116 -272 119 -270
rect 121 -272 124 -270
rect 116 -274 124 -272
rect 126 -267 134 -264
rect 126 -269 129 -267
rect 131 -269 134 -267
rect 126 -271 134 -269
rect 136 -259 144 -257
rect 136 -261 139 -259
rect 141 -261 144 -259
rect 136 -271 144 -261
rect 146 -259 153 -257
rect 146 -261 149 -259
rect 151 -261 153 -259
rect 146 -266 153 -261
rect 159 -264 164 -257
rect 146 -268 149 -266
rect 151 -268 153 -266
rect 146 -271 153 -268
rect 157 -266 164 -264
rect 157 -268 159 -266
rect 161 -268 164 -266
rect 157 -270 164 -268
rect 126 -274 131 -271
rect 116 -277 121 -274
rect 159 -277 164 -270
rect 166 -277 171 -257
rect 173 -263 180 -257
rect 173 -273 182 -263
rect 173 -275 176 -273
rect 178 -275 182 -273
rect 173 -277 182 -275
rect 184 -266 191 -263
rect 184 -268 187 -266
rect 189 -268 191 -266
rect 207 -264 214 -262
rect 207 -266 209 -264
rect 211 -266 214 -264
rect 207 -268 214 -266
rect 216 -264 224 -262
rect 216 -266 219 -264
rect 221 -266 224 -264
rect 216 -268 224 -266
rect 226 -264 234 -262
rect 226 -266 229 -264
rect 231 -266 234 -264
rect 226 -268 234 -266
rect 236 -264 243 -262
rect 270 -264 275 -257
rect 236 -266 239 -264
rect 241 -266 243 -264
rect 236 -268 243 -266
rect 248 -266 255 -264
rect 248 -268 250 -266
rect 252 -268 255 -266
rect 184 -270 191 -268
rect 184 -277 189 -270
rect 248 -270 255 -268
rect 250 -277 255 -270
rect 257 -270 265 -264
rect 257 -272 260 -270
rect 262 -272 265 -270
rect 257 -274 265 -272
rect 267 -267 275 -264
rect 267 -269 270 -267
rect 272 -269 275 -267
rect 267 -271 275 -269
rect 277 -259 285 -257
rect 277 -261 280 -259
rect 282 -261 285 -259
rect 277 -271 285 -261
rect 287 -259 294 -257
rect 287 -261 290 -259
rect 292 -261 294 -259
rect 287 -266 294 -261
rect 300 -264 305 -257
rect 287 -268 290 -266
rect 292 -268 294 -266
rect 287 -271 294 -268
rect 298 -266 305 -264
rect 298 -268 300 -266
rect 302 -268 305 -266
rect 298 -270 305 -268
rect 267 -274 272 -271
rect 257 -277 262 -274
rect 300 -277 305 -270
rect 307 -277 312 -257
rect 314 -263 321 -257
rect 314 -273 323 -263
rect 314 -275 317 -273
rect 319 -275 323 -273
rect 314 -277 323 -275
rect 325 -266 332 -263
rect 370 -264 375 -257
rect 325 -268 328 -266
rect 330 -268 332 -266
rect 325 -270 332 -268
rect 348 -266 355 -264
rect 348 -268 350 -266
rect 352 -268 355 -266
rect 348 -270 355 -268
rect 325 -277 330 -270
rect 350 -277 355 -270
rect 357 -270 365 -264
rect 357 -272 360 -270
rect 362 -272 365 -270
rect 357 -274 365 -272
rect 367 -267 375 -264
rect 367 -269 370 -267
rect 372 -269 375 -267
rect 367 -271 375 -269
rect 377 -259 385 -257
rect 377 -261 380 -259
rect 382 -261 385 -259
rect 377 -271 385 -261
rect 387 -259 394 -257
rect 387 -261 390 -259
rect 392 -261 394 -259
rect 387 -266 394 -261
rect 400 -264 405 -257
rect 387 -268 390 -266
rect 392 -268 394 -266
rect 387 -271 394 -268
rect 398 -266 405 -264
rect 398 -268 400 -266
rect 402 -268 405 -266
rect 398 -270 405 -268
rect 367 -274 372 -271
rect 357 -277 362 -274
rect 400 -277 405 -270
rect 407 -277 412 -257
rect 414 -263 421 -257
rect 414 -273 423 -263
rect 414 -275 417 -273
rect 419 -275 423 -273
rect 414 -277 423 -275
rect 425 -266 432 -263
rect 425 -268 428 -266
rect 430 -268 432 -266
rect 448 -264 455 -262
rect 448 -266 450 -264
rect 452 -266 455 -264
rect 448 -268 455 -266
rect 457 -264 465 -262
rect 457 -266 460 -264
rect 462 -266 465 -264
rect 457 -268 465 -266
rect 467 -264 475 -262
rect 467 -266 470 -264
rect 472 -266 475 -264
rect 467 -268 475 -266
rect 477 -264 484 -262
rect 477 -266 480 -264
rect 482 -266 484 -264
rect 477 -268 484 -266
rect 425 -270 432 -268
rect 425 -277 430 -270
<< pdif >>
rect 9 49 14 55
rect 7 47 14 49
rect 7 45 9 47
rect 11 45 14 47
rect 7 43 14 45
rect 16 53 22 55
rect 16 47 24 53
rect 16 45 19 47
rect 21 45 24 47
rect 16 43 24 45
rect 26 47 34 53
rect 26 45 29 47
rect 31 45 34 47
rect 26 43 34 45
rect 36 51 43 53
rect 36 49 39 51
rect 41 49 43 51
rect 53 49 58 55
rect 36 43 43 49
rect 51 47 58 49
rect 51 45 53 47
rect 55 45 58 47
rect 51 43 58 45
rect 60 53 66 55
rect 60 47 68 53
rect 60 45 63 47
rect 65 45 68 47
rect 60 43 68 45
rect 70 47 78 53
rect 70 45 73 47
rect 75 45 78 47
rect 70 43 78 45
rect 80 51 87 53
rect 80 49 83 51
rect 85 49 87 51
rect 97 49 102 55
rect 80 43 87 49
rect 95 47 102 49
rect 95 45 97 47
rect 99 45 102 47
rect 95 43 102 45
rect 104 53 110 55
rect 104 47 112 53
rect 104 45 107 47
rect 109 45 112 47
rect 104 43 112 45
rect 114 47 122 53
rect 114 45 117 47
rect 119 45 122 47
rect 114 43 122 45
rect 124 51 131 53
rect 124 49 127 51
rect 129 49 131 51
rect 141 49 146 55
rect 124 43 131 49
rect 139 47 146 49
rect 139 45 141 47
rect 143 45 146 47
rect 139 43 146 45
rect 148 53 154 55
rect 148 47 156 53
rect 148 45 151 47
rect 153 45 156 47
rect 148 43 156 45
rect 158 47 166 53
rect 158 45 161 47
rect 163 45 166 47
rect 158 43 166 45
rect 168 51 175 53
rect 168 49 171 51
rect 173 49 175 51
rect 185 49 190 55
rect 168 43 175 49
rect 183 47 190 49
rect 183 45 185 47
rect 187 45 190 47
rect 183 43 190 45
rect 192 53 198 55
rect 192 47 200 53
rect 192 45 195 47
rect 197 45 200 47
rect 192 43 200 45
rect 202 47 210 53
rect 202 45 205 47
rect 207 45 210 47
rect 202 43 210 45
rect 212 51 219 53
rect 212 49 215 51
rect 217 49 219 51
rect 229 49 234 55
rect 212 43 219 49
rect 227 47 234 49
rect 227 45 229 47
rect 231 45 234 47
rect 227 43 234 45
rect 236 53 242 55
rect 236 47 244 53
rect 236 45 239 47
rect 241 45 244 47
rect 236 43 244 45
rect 246 47 254 53
rect 246 45 249 47
rect 251 45 254 47
rect 246 43 254 45
rect 256 51 263 53
rect 256 49 259 51
rect 261 49 263 51
rect 273 49 278 55
rect 256 43 263 49
rect 271 47 278 49
rect 271 45 273 47
rect 275 45 278 47
rect 271 43 278 45
rect 280 53 286 55
rect 280 47 288 53
rect 280 45 283 47
rect 285 45 288 47
rect 280 43 288 45
rect 290 47 298 53
rect 290 45 293 47
rect 295 45 298 47
rect 290 43 298 45
rect 300 51 307 53
rect 300 49 303 51
rect 305 49 307 51
rect 317 49 322 55
rect 300 43 307 49
rect 315 47 322 49
rect 315 45 317 47
rect 319 45 322 47
rect 315 43 322 45
rect 324 53 330 55
rect 324 47 332 53
rect 324 45 327 47
rect 329 45 332 47
rect 324 43 332 45
rect 334 47 342 53
rect 334 45 337 47
rect 339 45 342 47
rect 334 43 342 45
rect 344 51 351 53
rect 344 49 347 51
rect 349 49 351 51
rect 361 49 366 55
rect 344 43 351 49
rect 359 47 366 49
rect 359 45 361 47
rect 363 45 366 47
rect 359 43 366 45
rect 368 53 374 55
rect 368 47 376 53
rect 368 45 371 47
rect 373 45 376 47
rect 368 43 376 45
rect 378 47 386 53
rect 378 45 381 47
rect 383 45 386 47
rect 378 43 386 45
rect 388 51 395 53
rect 388 49 391 51
rect 393 49 395 51
rect 405 49 410 55
rect 388 43 395 49
rect 403 47 410 49
rect 403 45 405 47
rect 407 45 410 47
rect 403 43 410 45
rect 412 53 418 55
rect 412 47 420 53
rect 412 45 415 47
rect 417 45 420 47
rect 412 43 420 45
rect 422 47 430 53
rect 422 45 425 47
rect 427 45 430 47
rect 422 43 430 45
rect 432 51 439 53
rect 432 49 435 51
rect 437 49 439 51
rect 449 49 454 55
rect 432 43 439 49
rect 447 47 454 49
rect 447 45 449 47
rect 451 45 454 47
rect 447 43 454 45
rect 456 53 462 55
rect 456 47 464 53
rect 456 45 459 47
rect 461 45 464 47
rect 456 43 464 45
rect 466 47 474 53
rect 466 45 469 47
rect 471 45 474 47
rect 466 43 474 45
rect 476 51 483 53
rect 476 49 479 51
rect 481 49 483 51
rect 493 49 498 55
rect 476 43 483 49
rect 491 47 498 49
rect 491 45 493 47
rect 495 45 498 47
rect 491 43 498 45
rect 500 53 506 55
rect 500 47 508 53
rect 500 45 503 47
rect 505 45 508 47
rect 500 43 508 45
rect 510 47 518 53
rect 510 45 513 47
rect 515 45 518 47
rect 510 43 518 45
rect 520 51 527 53
rect 520 49 523 51
rect 525 49 527 51
rect 537 49 542 55
rect 520 43 527 49
rect 535 47 542 49
rect 535 45 537 47
rect 539 45 542 47
rect 535 43 542 45
rect 544 53 550 55
rect 544 47 552 53
rect 544 45 547 47
rect 549 45 552 47
rect 544 43 552 45
rect 554 47 562 53
rect 554 45 557 47
rect 559 45 562 47
rect 554 43 562 45
rect 564 51 571 53
rect 564 49 567 51
rect 569 49 571 51
rect 581 49 586 55
rect 564 43 571 49
rect 579 47 586 49
rect 579 45 581 47
rect 583 45 586 47
rect 579 43 586 45
rect 588 53 594 55
rect 588 47 596 53
rect 588 45 591 47
rect 593 45 596 47
rect 588 43 596 45
rect 598 47 606 53
rect 598 45 601 47
rect 603 45 606 47
rect 598 43 606 45
rect 608 51 615 53
rect 608 49 611 51
rect 613 49 615 51
rect 625 49 630 55
rect 608 43 615 49
rect 623 47 630 49
rect 623 45 625 47
rect 627 45 630 47
rect 623 43 630 45
rect 632 53 638 55
rect 632 47 640 53
rect 632 45 635 47
rect 637 45 640 47
rect 632 43 640 45
rect 642 47 650 53
rect 642 45 645 47
rect 647 45 650 47
rect 642 43 650 45
rect 652 51 659 53
rect 652 49 655 51
rect 657 49 659 51
rect 669 49 674 55
rect 652 43 659 49
rect 667 47 674 49
rect 667 45 669 47
rect 671 45 674 47
rect 667 43 674 45
rect 676 53 682 55
rect 676 47 684 53
rect 676 45 679 47
rect 681 45 684 47
rect 676 43 684 45
rect 686 47 694 53
rect 686 45 689 47
rect 691 45 694 47
rect 686 43 694 45
rect 696 51 703 53
rect 696 49 699 51
rect 701 49 703 51
rect 696 43 703 49
rect 15 -35 22 -33
rect 15 -37 17 -35
rect 19 -37 22 -35
rect 15 -42 22 -37
rect 15 -44 17 -42
rect 19 -44 22 -42
rect 15 -46 22 -44
rect 17 -61 22 -46
rect 24 -50 32 -33
rect 24 -52 27 -50
rect 29 -52 32 -50
rect 24 -57 32 -52
rect 24 -59 27 -57
rect 29 -59 32 -57
rect 24 -61 32 -59
rect 34 -42 42 -33
rect 34 -44 37 -42
rect 39 -44 42 -42
rect 34 -49 42 -44
rect 34 -51 37 -49
rect 39 -51 42 -49
rect 34 -61 42 -51
rect 44 -50 60 -33
rect 44 -52 49 -50
rect 51 -52 60 -50
rect 44 -57 60 -52
rect 44 -59 49 -57
rect 51 -58 60 -57
rect 62 -58 67 -33
rect 69 -36 74 -33
rect 104 -35 111 -33
rect 69 -38 77 -36
rect 69 -40 72 -38
rect 74 -40 77 -38
rect 69 -49 77 -40
rect 79 -49 90 -36
rect 69 -58 74 -49
rect 81 -57 90 -49
rect 51 -59 58 -58
rect 44 -61 58 -59
rect 81 -59 84 -57
rect 86 -59 90 -57
rect 81 -61 90 -59
rect 92 -38 99 -36
rect 92 -40 95 -38
rect 97 -40 99 -38
rect 92 -45 99 -40
rect 92 -47 95 -45
rect 97 -47 99 -45
rect 104 -37 106 -35
rect 108 -37 111 -35
rect 104 -42 111 -37
rect 104 -44 106 -42
rect 108 -44 111 -42
rect 104 -46 111 -44
rect 92 -49 99 -47
rect 92 -61 97 -49
rect 106 -61 111 -46
rect 113 -50 121 -33
rect 113 -52 116 -50
rect 118 -52 121 -50
rect 113 -57 121 -52
rect 113 -59 116 -57
rect 118 -59 121 -57
rect 113 -61 121 -59
rect 123 -42 131 -33
rect 123 -44 126 -42
rect 128 -44 131 -42
rect 123 -49 131 -44
rect 123 -51 126 -49
rect 128 -51 131 -49
rect 123 -61 131 -51
rect 133 -50 149 -33
rect 133 -52 138 -50
rect 140 -52 149 -50
rect 133 -57 149 -52
rect 133 -59 138 -57
rect 140 -58 149 -57
rect 151 -58 156 -33
rect 158 -36 163 -33
rect 158 -38 166 -36
rect 158 -40 161 -38
rect 163 -40 166 -38
rect 158 -49 166 -40
rect 168 -49 179 -36
rect 158 -58 163 -49
rect 170 -57 179 -49
rect 140 -59 147 -58
rect 133 -61 147 -59
rect 170 -59 173 -57
rect 175 -59 179 -57
rect 170 -61 179 -59
rect 181 -38 188 -36
rect 181 -40 184 -38
rect 186 -40 188 -38
rect 181 -45 188 -40
rect 233 -35 240 -33
rect 233 -37 235 -35
rect 237 -37 240 -35
rect 211 -43 219 -40
rect 181 -47 184 -45
rect 186 -47 188 -45
rect 181 -49 188 -47
rect 194 -48 199 -43
rect 181 -61 186 -49
rect 192 -50 199 -48
rect 192 -52 194 -50
rect 196 -52 199 -50
rect 192 -54 199 -52
rect 194 -61 199 -54
rect 201 -61 206 -43
rect 208 -52 219 -43
rect 221 -46 226 -40
rect 233 -42 240 -37
rect 233 -44 235 -42
rect 237 -44 240 -42
rect 233 -46 240 -44
rect 221 -48 228 -46
rect 221 -50 224 -48
rect 226 -50 228 -48
rect 221 -52 228 -50
rect 208 -57 217 -52
rect 208 -59 212 -57
rect 214 -59 217 -57
rect 208 -61 217 -59
rect 235 -61 240 -46
rect 242 -50 250 -33
rect 242 -52 245 -50
rect 247 -52 250 -50
rect 242 -57 250 -52
rect 242 -59 245 -57
rect 247 -59 250 -57
rect 242 -61 250 -59
rect 252 -42 260 -33
rect 252 -44 255 -42
rect 257 -44 260 -42
rect 252 -49 260 -44
rect 252 -51 255 -49
rect 257 -51 260 -49
rect 252 -61 260 -51
rect 262 -50 278 -33
rect 262 -52 267 -50
rect 269 -52 278 -50
rect 262 -57 278 -52
rect 262 -59 267 -57
rect 269 -58 278 -57
rect 280 -58 285 -33
rect 287 -36 292 -33
rect 322 -35 329 -33
rect 287 -38 295 -36
rect 287 -40 290 -38
rect 292 -40 295 -38
rect 287 -49 295 -40
rect 297 -49 308 -36
rect 287 -58 292 -49
rect 299 -57 308 -49
rect 269 -59 276 -58
rect 262 -61 276 -59
rect 299 -59 302 -57
rect 304 -59 308 -57
rect 299 -61 308 -59
rect 310 -38 317 -36
rect 310 -40 313 -38
rect 315 -40 317 -38
rect 310 -45 317 -40
rect 310 -47 313 -45
rect 315 -47 317 -45
rect 322 -37 324 -35
rect 326 -37 329 -35
rect 322 -42 329 -37
rect 322 -44 324 -42
rect 326 -44 329 -42
rect 322 -46 329 -44
rect 310 -49 317 -47
rect 310 -61 315 -49
rect 324 -61 329 -46
rect 331 -50 339 -33
rect 331 -52 334 -50
rect 336 -52 339 -50
rect 331 -57 339 -52
rect 331 -59 334 -57
rect 336 -59 339 -57
rect 331 -61 339 -59
rect 341 -42 349 -33
rect 341 -44 344 -42
rect 346 -44 349 -42
rect 341 -49 349 -44
rect 341 -51 344 -49
rect 346 -51 349 -49
rect 341 -61 349 -51
rect 351 -50 367 -33
rect 351 -52 356 -50
rect 358 -52 367 -50
rect 351 -57 367 -52
rect 351 -59 356 -57
rect 358 -58 367 -57
rect 369 -58 374 -33
rect 376 -36 381 -33
rect 491 -35 498 -33
rect 376 -38 384 -36
rect 376 -40 379 -38
rect 381 -40 384 -38
rect 376 -49 384 -40
rect 386 -49 397 -36
rect 376 -58 381 -49
rect 388 -57 397 -49
rect 358 -59 365 -58
rect 351 -61 365 -59
rect 388 -59 391 -57
rect 393 -59 397 -57
rect 388 -61 397 -59
rect 399 -38 406 -36
rect 399 -40 402 -38
rect 404 -40 406 -38
rect 399 -45 406 -40
rect 399 -47 402 -45
rect 404 -47 406 -45
rect 491 -37 493 -35
rect 495 -37 498 -35
rect 491 -42 498 -37
rect 491 -44 493 -42
rect 495 -44 498 -42
rect 491 -46 498 -44
rect 399 -49 406 -47
rect 399 -61 404 -49
rect 493 -61 498 -46
rect 500 -50 508 -33
rect 500 -52 503 -50
rect 505 -52 508 -50
rect 500 -57 508 -52
rect 500 -59 503 -57
rect 505 -59 508 -57
rect 500 -61 508 -59
rect 510 -42 518 -33
rect 510 -44 513 -42
rect 515 -44 518 -42
rect 510 -49 518 -44
rect 510 -51 513 -49
rect 515 -51 518 -49
rect 510 -61 518 -51
rect 520 -50 536 -33
rect 520 -52 525 -50
rect 527 -52 536 -50
rect 520 -57 536 -52
rect 520 -59 525 -57
rect 527 -58 536 -57
rect 538 -58 543 -33
rect 545 -36 550 -33
rect 580 -35 587 -33
rect 545 -38 553 -36
rect 545 -40 548 -38
rect 550 -40 553 -38
rect 545 -49 553 -40
rect 555 -49 566 -36
rect 545 -58 550 -49
rect 557 -57 566 -49
rect 527 -59 534 -58
rect 520 -61 534 -59
rect 557 -59 560 -57
rect 562 -59 566 -57
rect 557 -61 566 -59
rect 568 -38 575 -36
rect 568 -40 571 -38
rect 573 -40 575 -38
rect 568 -45 575 -40
rect 568 -47 571 -45
rect 573 -47 575 -45
rect 580 -37 582 -35
rect 584 -37 587 -35
rect 580 -42 587 -37
rect 580 -44 582 -42
rect 584 -44 587 -42
rect 580 -46 587 -44
rect 568 -49 575 -47
rect 568 -61 573 -49
rect 582 -61 587 -46
rect 589 -50 597 -33
rect 589 -52 592 -50
rect 594 -52 597 -50
rect 589 -57 597 -52
rect 589 -59 592 -57
rect 594 -59 597 -57
rect 589 -61 597 -59
rect 599 -42 607 -33
rect 599 -44 602 -42
rect 604 -44 607 -42
rect 599 -49 607 -44
rect 599 -51 602 -49
rect 604 -51 607 -49
rect 599 -61 607 -51
rect 609 -50 625 -33
rect 609 -52 614 -50
rect 616 -52 625 -50
rect 609 -57 625 -52
rect 609 -59 614 -57
rect 616 -58 625 -57
rect 627 -58 632 -33
rect 634 -36 639 -33
rect 634 -38 642 -36
rect 634 -40 637 -38
rect 639 -40 642 -38
rect 634 -49 642 -40
rect 644 -49 655 -36
rect 634 -58 639 -49
rect 646 -57 655 -49
rect 616 -59 623 -58
rect 609 -61 623 -59
rect 646 -59 649 -57
rect 651 -59 655 -57
rect 646 -61 655 -59
rect 657 -38 664 -36
rect 657 -40 660 -38
rect 662 -40 664 -38
rect 657 -45 664 -40
rect 657 -47 660 -45
rect 662 -47 664 -45
rect 657 -49 664 -47
rect 657 -61 662 -49
rect 9 -85 14 -73
rect 7 -87 14 -85
rect 7 -89 9 -87
rect 11 -89 14 -87
rect 7 -94 14 -89
rect 7 -96 9 -94
rect 11 -96 14 -94
rect 7 -98 14 -96
rect 16 -75 25 -73
rect 16 -77 20 -75
rect 22 -77 25 -75
rect 48 -75 62 -73
rect 48 -76 55 -75
rect 16 -85 25 -77
rect 32 -85 37 -76
rect 16 -98 27 -85
rect 29 -94 37 -85
rect 29 -96 32 -94
rect 34 -96 37 -94
rect 29 -98 37 -96
rect 32 -101 37 -98
rect 39 -101 44 -76
rect 46 -77 55 -76
rect 57 -77 62 -75
rect 46 -82 62 -77
rect 46 -84 55 -82
rect 57 -84 62 -82
rect 46 -101 62 -84
rect 64 -83 72 -73
rect 64 -85 67 -83
rect 69 -85 72 -83
rect 64 -90 72 -85
rect 64 -92 67 -90
rect 69 -92 72 -90
rect 64 -101 72 -92
rect 74 -75 82 -73
rect 74 -77 77 -75
rect 79 -77 82 -75
rect 74 -82 82 -77
rect 74 -84 77 -82
rect 79 -84 82 -82
rect 74 -101 82 -84
rect 84 -88 89 -73
rect 98 -85 103 -73
rect 96 -87 103 -85
rect 84 -90 91 -88
rect 84 -92 87 -90
rect 89 -92 91 -90
rect 84 -97 91 -92
rect 84 -99 87 -97
rect 89 -99 91 -97
rect 96 -89 98 -87
rect 100 -89 103 -87
rect 96 -94 103 -89
rect 96 -96 98 -94
rect 100 -96 103 -94
rect 96 -98 103 -96
rect 105 -75 114 -73
rect 105 -77 109 -75
rect 111 -77 114 -75
rect 137 -75 151 -73
rect 137 -76 144 -75
rect 105 -85 114 -77
rect 121 -85 126 -76
rect 105 -98 116 -85
rect 118 -94 126 -85
rect 118 -96 121 -94
rect 123 -96 126 -94
rect 118 -98 126 -96
rect 84 -101 91 -99
rect 121 -101 126 -98
rect 128 -101 133 -76
rect 135 -77 144 -76
rect 146 -77 151 -75
rect 135 -82 151 -77
rect 135 -84 144 -82
rect 146 -84 151 -82
rect 135 -101 151 -84
rect 153 -83 161 -73
rect 153 -85 156 -83
rect 158 -85 161 -83
rect 153 -90 161 -85
rect 153 -92 156 -90
rect 158 -92 161 -90
rect 153 -101 161 -92
rect 163 -75 171 -73
rect 163 -77 166 -75
rect 168 -77 171 -75
rect 163 -82 171 -77
rect 163 -84 166 -82
rect 168 -84 171 -82
rect 163 -101 171 -84
rect 173 -88 178 -73
rect 196 -75 205 -73
rect 196 -77 199 -75
rect 201 -77 205 -75
rect 196 -82 205 -77
rect 185 -84 192 -82
rect 185 -86 187 -84
rect 189 -86 192 -84
rect 185 -88 192 -86
rect 173 -90 180 -88
rect 173 -92 176 -90
rect 178 -92 180 -90
rect 173 -97 180 -92
rect 187 -94 192 -88
rect 194 -91 205 -82
rect 207 -91 212 -73
rect 214 -80 219 -73
rect 214 -82 221 -80
rect 214 -84 217 -82
rect 219 -84 221 -82
rect 214 -86 221 -84
rect 227 -85 232 -73
rect 214 -91 219 -86
rect 225 -87 232 -85
rect 225 -89 227 -87
rect 229 -89 232 -87
rect 194 -94 202 -91
rect 173 -99 176 -97
rect 178 -99 180 -97
rect 173 -101 180 -99
rect 225 -94 232 -89
rect 225 -96 227 -94
rect 229 -96 232 -94
rect 225 -98 232 -96
rect 234 -75 243 -73
rect 234 -77 238 -75
rect 240 -77 243 -75
rect 266 -75 280 -73
rect 266 -76 273 -75
rect 234 -85 243 -77
rect 250 -85 255 -76
rect 234 -98 245 -85
rect 247 -94 255 -85
rect 247 -96 250 -94
rect 252 -96 255 -94
rect 247 -98 255 -96
rect 250 -101 255 -98
rect 257 -101 262 -76
rect 264 -77 273 -76
rect 275 -77 280 -75
rect 264 -82 280 -77
rect 264 -84 273 -82
rect 275 -84 280 -82
rect 264 -101 280 -84
rect 282 -83 290 -73
rect 282 -85 285 -83
rect 287 -85 290 -83
rect 282 -90 290 -85
rect 282 -92 285 -90
rect 287 -92 290 -90
rect 282 -101 290 -92
rect 292 -75 300 -73
rect 292 -77 295 -75
rect 297 -77 300 -75
rect 292 -82 300 -77
rect 292 -84 295 -82
rect 297 -84 300 -82
rect 292 -101 300 -84
rect 302 -88 307 -73
rect 316 -85 321 -73
rect 314 -87 321 -85
rect 302 -90 309 -88
rect 302 -92 305 -90
rect 307 -92 309 -90
rect 302 -97 309 -92
rect 302 -99 305 -97
rect 307 -99 309 -97
rect 314 -89 316 -87
rect 318 -89 321 -87
rect 314 -94 321 -89
rect 314 -96 316 -94
rect 318 -96 321 -94
rect 314 -98 321 -96
rect 323 -75 332 -73
rect 323 -77 327 -75
rect 329 -77 332 -75
rect 355 -75 369 -73
rect 355 -76 362 -75
rect 323 -85 332 -77
rect 339 -85 344 -76
rect 323 -98 334 -85
rect 336 -94 344 -85
rect 336 -96 339 -94
rect 341 -96 344 -94
rect 336 -98 344 -96
rect 302 -101 309 -99
rect 339 -101 344 -98
rect 346 -101 351 -76
rect 353 -77 362 -76
rect 364 -77 369 -75
rect 353 -82 369 -77
rect 353 -84 362 -82
rect 364 -84 369 -82
rect 353 -101 369 -84
rect 371 -83 379 -73
rect 371 -85 374 -83
rect 376 -85 379 -83
rect 371 -90 379 -85
rect 371 -92 374 -90
rect 376 -92 379 -90
rect 371 -101 379 -92
rect 381 -75 389 -73
rect 381 -77 384 -75
rect 386 -77 389 -75
rect 381 -82 389 -77
rect 381 -84 384 -82
rect 386 -84 389 -82
rect 381 -101 389 -84
rect 391 -88 396 -73
rect 414 -75 423 -73
rect 414 -77 417 -75
rect 419 -77 423 -75
rect 414 -82 423 -77
rect 403 -84 410 -82
rect 403 -86 405 -84
rect 407 -86 410 -84
rect 403 -88 410 -86
rect 391 -90 398 -88
rect 391 -92 394 -90
rect 396 -92 398 -90
rect 391 -97 398 -92
rect 405 -94 410 -88
rect 412 -91 423 -82
rect 425 -91 430 -73
rect 432 -80 437 -73
rect 432 -82 439 -80
rect 432 -84 435 -82
rect 437 -84 439 -82
rect 432 -86 439 -84
rect 445 -85 450 -73
rect 432 -91 437 -86
rect 443 -87 450 -85
rect 443 -89 445 -87
rect 447 -89 450 -87
rect 412 -94 420 -91
rect 391 -99 394 -97
rect 396 -99 398 -97
rect 391 -101 398 -99
rect 443 -94 450 -89
rect 443 -96 445 -94
rect 447 -96 450 -94
rect 443 -98 450 -96
rect 452 -75 461 -73
rect 452 -77 456 -75
rect 458 -77 461 -75
rect 484 -75 498 -73
rect 484 -76 491 -75
rect 452 -85 461 -77
rect 468 -85 473 -76
rect 452 -98 463 -85
rect 465 -94 473 -85
rect 465 -96 468 -94
rect 470 -96 473 -94
rect 465 -98 473 -96
rect 468 -101 473 -98
rect 475 -101 480 -76
rect 482 -77 491 -76
rect 493 -77 498 -75
rect 482 -82 498 -77
rect 482 -84 491 -82
rect 493 -84 498 -82
rect 482 -101 498 -84
rect 500 -83 508 -73
rect 500 -85 503 -83
rect 505 -85 508 -83
rect 500 -90 508 -85
rect 500 -92 503 -90
rect 505 -92 508 -90
rect 500 -101 508 -92
rect 510 -75 518 -73
rect 510 -77 513 -75
rect 515 -77 518 -75
rect 510 -82 518 -77
rect 510 -84 513 -82
rect 515 -84 518 -82
rect 510 -101 518 -84
rect 520 -88 525 -73
rect 534 -85 539 -73
rect 532 -87 539 -85
rect 520 -90 527 -88
rect 520 -92 523 -90
rect 525 -92 527 -90
rect 520 -97 527 -92
rect 520 -99 523 -97
rect 525 -99 527 -97
rect 532 -89 534 -87
rect 536 -89 539 -87
rect 532 -94 539 -89
rect 532 -96 534 -94
rect 536 -96 539 -94
rect 532 -98 539 -96
rect 541 -75 550 -73
rect 541 -77 545 -75
rect 547 -77 550 -75
rect 573 -75 587 -73
rect 573 -76 580 -75
rect 541 -85 550 -77
rect 557 -85 562 -76
rect 541 -98 552 -85
rect 554 -94 562 -85
rect 554 -96 557 -94
rect 559 -96 562 -94
rect 554 -98 562 -96
rect 520 -101 527 -99
rect 557 -101 562 -98
rect 564 -101 569 -76
rect 571 -77 580 -76
rect 582 -77 587 -75
rect 571 -82 587 -77
rect 571 -84 580 -82
rect 582 -84 587 -82
rect 571 -101 587 -84
rect 589 -83 597 -73
rect 589 -85 592 -83
rect 594 -85 597 -83
rect 589 -90 597 -85
rect 589 -92 592 -90
rect 594 -92 597 -90
rect 589 -101 597 -92
rect 599 -75 607 -73
rect 599 -77 602 -75
rect 604 -77 607 -75
rect 599 -82 607 -77
rect 599 -84 602 -82
rect 604 -84 607 -82
rect 599 -101 607 -84
rect 609 -88 614 -73
rect 632 -75 641 -73
rect 632 -77 635 -75
rect 637 -77 641 -75
rect 632 -82 641 -77
rect 621 -84 628 -82
rect 621 -86 623 -84
rect 625 -86 628 -84
rect 621 -88 628 -86
rect 609 -90 616 -88
rect 609 -92 612 -90
rect 614 -92 616 -90
rect 609 -97 616 -92
rect 623 -94 628 -88
rect 630 -91 641 -82
rect 643 -91 648 -73
rect 650 -80 655 -73
rect 650 -82 657 -80
rect 650 -84 653 -82
rect 655 -84 657 -82
rect 650 -86 657 -84
rect 650 -91 655 -86
rect 630 -94 638 -91
rect 609 -99 612 -97
rect 614 -99 616 -97
rect 609 -101 616 -99
rect 284 -179 291 -177
rect 284 -181 286 -179
rect 288 -181 291 -179
rect 251 -187 259 -184
rect 234 -192 239 -187
rect 232 -194 239 -192
rect 232 -196 234 -194
rect 236 -196 239 -194
rect 232 -198 239 -196
rect 234 -205 239 -198
rect 241 -205 246 -187
rect 248 -196 259 -187
rect 261 -190 266 -184
rect 284 -186 291 -181
rect 284 -188 286 -186
rect 288 -188 291 -186
rect 284 -190 291 -188
rect 261 -192 268 -190
rect 261 -194 264 -192
rect 266 -194 268 -192
rect 261 -196 268 -194
rect 248 -201 257 -196
rect 248 -203 252 -201
rect 254 -203 257 -201
rect 248 -205 257 -203
rect 286 -205 291 -190
rect 293 -194 301 -177
rect 293 -196 296 -194
rect 298 -196 301 -194
rect 293 -201 301 -196
rect 293 -203 296 -201
rect 298 -203 301 -201
rect 293 -205 301 -203
rect 303 -186 311 -177
rect 303 -188 306 -186
rect 308 -188 311 -186
rect 303 -193 311 -188
rect 303 -195 306 -193
rect 308 -195 311 -193
rect 303 -205 311 -195
rect 313 -194 329 -177
rect 313 -196 318 -194
rect 320 -196 329 -194
rect 313 -201 329 -196
rect 313 -203 318 -201
rect 320 -202 329 -201
rect 331 -202 336 -177
rect 338 -180 343 -177
rect 384 -179 391 -177
rect 338 -182 346 -180
rect 338 -184 341 -182
rect 343 -184 346 -182
rect 338 -193 346 -184
rect 348 -193 359 -180
rect 338 -202 343 -193
rect 350 -201 359 -193
rect 320 -203 327 -202
rect 313 -205 327 -203
rect 350 -203 353 -201
rect 355 -203 359 -201
rect 350 -205 359 -203
rect 361 -182 368 -180
rect 361 -184 364 -182
rect 366 -184 368 -182
rect 361 -189 368 -184
rect 361 -191 364 -189
rect 366 -191 368 -189
rect 384 -181 386 -179
rect 388 -181 391 -179
rect 384 -186 391 -181
rect 384 -188 386 -186
rect 388 -188 391 -186
rect 384 -190 391 -188
rect 361 -193 368 -191
rect 361 -205 366 -193
rect 386 -205 391 -190
rect 393 -194 401 -177
rect 393 -196 396 -194
rect 398 -196 401 -194
rect 393 -201 401 -196
rect 393 -203 396 -201
rect 398 -203 401 -201
rect 393 -205 401 -203
rect 403 -186 411 -177
rect 403 -188 406 -186
rect 408 -188 411 -186
rect 403 -193 411 -188
rect 403 -195 406 -193
rect 408 -195 411 -193
rect 403 -205 411 -195
rect 413 -194 429 -177
rect 413 -196 418 -194
rect 420 -196 429 -194
rect 413 -201 429 -196
rect 413 -203 418 -201
rect 420 -202 429 -201
rect 431 -202 436 -177
rect 438 -180 443 -177
rect 438 -182 446 -180
rect 438 -184 441 -182
rect 443 -184 446 -182
rect 438 -193 446 -184
rect 448 -193 459 -180
rect 438 -202 443 -193
rect 450 -201 459 -193
rect 420 -203 427 -202
rect 413 -205 427 -203
rect 450 -203 453 -201
rect 455 -203 459 -201
rect 450 -205 459 -203
rect 461 -182 468 -180
rect 461 -184 464 -182
rect 466 -184 468 -182
rect 461 -189 468 -184
rect 528 -179 535 -177
rect 528 -181 530 -179
rect 532 -181 535 -179
rect 495 -187 503 -184
rect 461 -191 464 -189
rect 466 -191 468 -189
rect 461 -193 468 -191
rect 478 -192 483 -187
rect 461 -205 466 -193
rect 476 -194 483 -192
rect 476 -196 478 -194
rect 480 -196 483 -194
rect 476 -198 483 -196
rect 478 -205 483 -198
rect 485 -205 490 -187
rect 492 -196 503 -187
rect 505 -190 510 -184
rect 528 -186 535 -181
rect 528 -188 530 -186
rect 532 -188 535 -186
rect 528 -190 535 -188
rect 505 -192 512 -190
rect 505 -194 508 -192
rect 510 -194 512 -192
rect 505 -196 512 -194
rect 492 -201 501 -196
rect 492 -203 496 -201
rect 498 -203 501 -201
rect 492 -205 501 -203
rect 530 -205 535 -190
rect 537 -194 545 -177
rect 537 -196 540 -194
rect 542 -196 545 -194
rect 537 -201 545 -196
rect 537 -203 540 -201
rect 542 -203 545 -201
rect 537 -205 545 -203
rect 547 -186 555 -177
rect 547 -188 550 -186
rect 552 -188 555 -186
rect 547 -193 555 -188
rect 547 -195 550 -193
rect 552 -195 555 -193
rect 547 -205 555 -195
rect 557 -194 573 -177
rect 557 -196 562 -194
rect 564 -196 573 -194
rect 557 -201 573 -196
rect 557 -203 562 -201
rect 564 -202 573 -201
rect 575 -202 580 -177
rect 582 -180 587 -177
rect 628 -179 635 -177
rect 582 -182 590 -180
rect 582 -184 585 -182
rect 587 -184 590 -182
rect 582 -193 590 -184
rect 592 -193 603 -180
rect 582 -202 587 -193
rect 594 -201 603 -193
rect 564 -203 571 -202
rect 557 -205 571 -203
rect 594 -203 597 -201
rect 599 -203 603 -201
rect 594 -205 603 -203
rect 605 -182 612 -180
rect 605 -184 608 -182
rect 610 -184 612 -182
rect 605 -189 612 -184
rect 605 -191 608 -189
rect 610 -191 612 -189
rect 628 -181 630 -179
rect 632 -181 635 -179
rect 628 -186 635 -181
rect 628 -188 630 -186
rect 632 -188 635 -186
rect 628 -190 635 -188
rect 605 -193 612 -191
rect 605 -205 610 -193
rect 630 -205 635 -190
rect 637 -194 645 -177
rect 637 -196 640 -194
rect 642 -196 645 -194
rect 637 -201 645 -196
rect 637 -203 640 -201
rect 642 -203 645 -201
rect 637 -205 645 -203
rect 647 -186 655 -177
rect 647 -188 650 -186
rect 652 -188 655 -186
rect 647 -193 655 -188
rect 647 -195 650 -193
rect 652 -195 655 -193
rect 647 -205 655 -195
rect 657 -194 673 -177
rect 657 -196 662 -194
rect 664 -196 673 -194
rect 657 -201 673 -196
rect 657 -203 662 -201
rect 664 -202 673 -201
rect 675 -202 680 -177
rect 682 -180 687 -177
rect 682 -182 690 -180
rect 682 -184 685 -182
rect 687 -184 690 -182
rect 682 -193 690 -184
rect 692 -193 703 -180
rect 682 -202 687 -193
rect 694 -201 703 -193
rect 664 -203 671 -202
rect 657 -205 671 -203
rect 694 -203 697 -201
rect 699 -203 703 -201
rect 694 -205 703 -203
rect 705 -182 712 -180
rect 705 -184 708 -182
rect 710 -184 712 -182
rect 705 -189 712 -184
rect 705 -191 708 -189
rect 710 -191 712 -189
rect 705 -193 712 -191
rect 705 -205 710 -193
rect 9 -229 14 -217
rect 7 -231 14 -229
rect 7 -233 9 -231
rect 11 -233 14 -231
rect 7 -238 14 -233
rect 7 -240 9 -238
rect 11 -240 14 -238
rect 7 -242 14 -240
rect 16 -219 25 -217
rect 16 -221 20 -219
rect 22 -221 25 -219
rect 48 -219 62 -217
rect 48 -220 55 -219
rect 16 -229 25 -221
rect 32 -229 37 -220
rect 16 -242 27 -229
rect 29 -238 37 -229
rect 29 -240 32 -238
rect 34 -240 37 -238
rect 29 -242 37 -240
rect 32 -245 37 -242
rect 39 -245 44 -220
rect 46 -221 55 -220
rect 57 -221 62 -219
rect 46 -226 62 -221
rect 46 -228 55 -226
rect 57 -228 62 -226
rect 46 -245 62 -228
rect 64 -227 72 -217
rect 64 -229 67 -227
rect 69 -229 72 -227
rect 64 -234 72 -229
rect 64 -236 67 -234
rect 69 -236 72 -234
rect 64 -245 72 -236
rect 74 -219 82 -217
rect 74 -221 77 -219
rect 79 -221 82 -219
rect 74 -226 82 -221
rect 74 -228 77 -226
rect 79 -228 82 -226
rect 74 -245 82 -228
rect 84 -232 89 -217
rect 109 -229 114 -217
rect 107 -231 114 -229
rect 84 -234 91 -232
rect 84 -236 87 -234
rect 89 -236 91 -234
rect 84 -241 91 -236
rect 84 -243 87 -241
rect 89 -243 91 -241
rect 107 -233 109 -231
rect 111 -233 114 -231
rect 107 -238 114 -233
rect 107 -240 109 -238
rect 111 -240 114 -238
rect 107 -242 114 -240
rect 116 -219 125 -217
rect 116 -221 120 -219
rect 122 -221 125 -219
rect 148 -219 162 -217
rect 148 -220 155 -219
rect 116 -229 125 -221
rect 132 -229 137 -220
rect 116 -242 127 -229
rect 129 -238 137 -229
rect 129 -240 132 -238
rect 134 -240 137 -238
rect 129 -242 137 -240
rect 84 -245 91 -243
rect 132 -245 137 -242
rect 139 -245 144 -220
rect 146 -221 155 -220
rect 157 -221 162 -219
rect 146 -226 162 -221
rect 146 -228 155 -226
rect 157 -228 162 -226
rect 146 -245 162 -228
rect 164 -227 172 -217
rect 164 -229 167 -227
rect 169 -229 172 -227
rect 164 -234 172 -229
rect 164 -236 167 -234
rect 169 -236 172 -234
rect 164 -245 172 -236
rect 174 -219 182 -217
rect 174 -221 177 -219
rect 179 -221 182 -219
rect 174 -226 182 -221
rect 174 -228 177 -226
rect 179 -228 182 -226
rect 174 -245 182 -228
rect 184 -232 189 -217
rect 218 -219 227 -217
rect 218 -221 221 -219
rect 223 -221 227 -219
rect 218 -226 227 -221
rect 207 -228 214 -226
rect 207 -230 209 -228
rect 211 -230 214 -228
rect 207 -232 214 -230
rect 184 -234 191 -232
rect 184 -236 187 -234
rect 189 -236 191 -234
rect 184 -241 191 -236
rect 209 -238 214 -232
rect 216 -235 227 -226
rect 229 -235 234 -217
rect 236 -224 241 -217
rect 236 -226 243 -224
rect 236 -228 239 -226
rect 241 -228 243 -226
rect 236 -230 243 -228
rect 250 -229 255 -217
rect 236 -235 241 -230
rect 248 -231 255 -229
rect 248 -233 250 -231
rect 252 -233 255 -231
rect 216 -238 224 -235
rect 184 -243 187 -241
rect 189 -243 191 -241
rect 184 -245 191 -243
rect 248 -238 255 -233
rect 248 -240 250 -238
rect 252 -240 255 -238
rect 248 -242 255 -240
rect 257 -219 266 -217
rect 257 -221 261 -219
rect 263 -221 266 -219
rect 289 -219 303 -217
rect 289 -220 296 -219
rect 257 -229 266 -221
rect 273 -229 278 -220
rect 257 -242 268 -229
rect 270 -238 278 -229
rect 270 -240 273 -238
rect 275 -240 278 -238
rect 270 -242 278 -240
rect 273 -245 278 -242
rect 280 -245 285 -220
rect 287 -221 296 -220
rect 298 -221 303 -219
rect 287 -226 303 -221
rect 287 -228 296 -226
rect 298 -228 303 -226
rect 287 -245 303 -228
rect 305 -227 313 -217
rect 305 -229 308 -227
rect 310 -229 313 -227
rect 305 -234 313 -229
rect 305 -236 308 -234
rect 310 -236 313 -234
rect 305 -245 313 -236
rect 315 -219 323 -217
rect 315 -221 318 -219
rect 320 -221 323 -219
rect 315 -226 323 -221
rect 315 -228 318 -226
rect 320 -228 323 -226
rect 315 -245 323 -228
rect 325 -232 330 -217
rect 350 -229 355 -217
rect 348 -231 355 -229
rect 325 -234 332 -232
rect 325 -236 328 -234
rect 330 -236 332 -234
rect 325 -241 332 -236
rect 325 -243 328 -241
rect 330 -243 332 -241
rect 348 -233 350 -231
rect 352 -233 355 -231
rect 348 -238 355 -233
rect 348 -240 350 -238
rect 352 -240 355 -238
rect 348 -242 355 -240
rect 357 -219 366 -217
rect 357 -221 361 -219
rect 363 -221 366 -219
rect 389 -219 403 -217
rect 389 -220 396 -219
rect 357 -229 366 -221
rect 373 -229 378 -220
rect 357 -242 368 -229
rect 370 -238 378 -229
rect 370 -240 373 -238
rect 375 -240 378 -238
rect 370 -242 378 -240
rect 325 -245 332 -243
rect 373 -245 378 -242
rect 380 -245 385 -220
rect 387 -221 396 -220
rect 398 -221 403 -219
rect 387 -226 403 -221
rect 387 -228 396 -226
rect 398 -228 403 -226
rect 387 -245 403 -228
rect 405 -227 413 -217
rect 405 -229 408 -227
rect 410 -229 413 -227
rect 405 -234 413 -229
rect 405 -236 408 -234
rect 410 -236 413 -234
rect 405 -245 413 -236
rect 415 -219 423 -217
rect 415 -221 418 -219
rect 420 -221 423 -219
rect 415 -226 423 -221
rect 415 -228 418 -226
rect 420 -228 423 -226
rect 415 -245 423 -228
rect 425 -232 430 -217
rect 459 -219 468 -217
rect 459 -221 462 -219
rect 464 -221 468 -219
rect 459 -226 468 -221
rect 448 -228 455 -226
rect 448 -230 450 -228
rect 452 -230 455 -228
rect 448 -232 455 -230
rect 425 -234 432 -232
rect 425 -236 428 -234
rect 430 -236 432 -234
rect 425 -241 432 -236
rect 450 -238 455 -232
rect 457 -235 468 -226
rect 470 -235 475 -217
rect 477 -224 482 -217
rect 477 -226 484 -224
rect 477 -228 480 -226
rect 482 -228 484 -226
rect 477 -230 484 -228
rect 477 -235 482 -230
rect 457 -238 465 -235
rect 425 -243 428 -241
rect 430 -243 432 -241
rect 425 -245 432 -243
<< alu1 >>
rect 39 142 307 143
rect 39 140 40 142
rect 42 140 84 142
rect 86 140 172 142
rect 174 140 304 142
rect 306 140 307 142
rect 39 139 307 140
rect 31 134 431 135
rect 31 132 32 134
rect 34 132 120 134
rect 122 132 252 134
rect 254 132 428 134
rect 430 132 431 134
rect 31 131 431 132
rect 127 126 571 127
rect 127 124 128 126
rect 130 124 216 126
rect 218 124 348 126
rect 350 124 568 126
rect 570 124 571 126
rect 127 123 571 124
rect 75 118 475 119
rect 75 116 76 118
rect 78 116 208 118
rect 210 116 384 118
rect 386 116 472 118
rect 474 116 475 118
rect 75 115 475 116
rect 258 110 615 111
rect 258 108 260 110
rect 262 108 392 110
rect 394 108 524 110
rect 526 108 612 110
rect 614 108 615 110
rect 258 107 615 108
rect 163 102 651 103
rect 163 100 164 102
rect 166 100 340 102
rect 342 100 516 102
rect 518 100 648 102
rect 650 100 651 102
rect 163 99 651 100
rect 435 94 707 95
rect 435 92 436 94
rect 438 92 480 94
rect 482 92 656 94
rect 658 92 700 94
rect 702 92 707 94
rect 435 91 707 92
rect 295 86 707 87
rect 295 84 296 86
rect 298 84 560 86
rect 562 84 604 86
rect 606 84 692 86
rect 694 84 707 86
rect 295 83 707 84
rect -22 74 738 77
rect -22 72 -19 74
rect -17 72 733 74
rect 735 72 738 74
rect -22 70 10 72
rect 12 70 24 72
rect 26 70 38 72
rect 40 70 54 72
rect 56 70 68 72
rect 70 70 82 72
rect 84 70 98 72
rect 100 70 112 72
rect 114 70 126 72
rect 128 70 142 72
rect 144 70 156 72
rect 158 70 170 72
rect 172 70 186 72
rect 188 70 200 72
rect 202 70 214 72
rect 216 70 230 72
rect 232 70 244 72
rect 246 70 258 72
rect 260 70 274 72
rect 276 70 288 72
rect 290 70 302 72
rect 304 70 318 72
rect 320 70 332 72
rect 334 70 346 72
rect 348 70 362 72
rect 364 70 376 72
rect 378 70 390 72
rect 392 70 406 72
rect 408 70 420 72
rect 422 70 434 72
rect 436 70 450 72
rect 452 70 464 72
rect 466 70 478 72
rect 480 70 494 72
rect 496 70 508 72
rect 510 70 522 72
rect 524 70 538 72
rect 540 70 552 72
rect 554 70 566 72
rect 568 70 582 72
rect 584 70 596 72
rect 598 70 610 72
rect 612 70 626 72
rect 628 70 640 72
rect 642 70 654 72
rect 656 70 670 72
rect 672 70 684 72
rect 686 70 698 72
rect 700 70 738 72
rect -22 69 738 70
rect 7 47 11 56
rect 7 45 9 47
rect 7 31 11 45
rect 22 63 35 64
rect 22 62 32 63
rect 22 60 26 62
rect 28 61 32 62
rect 34 61 35 63
rect 28 60 35 61
rect 22 58 35 60
rect 22 51 28 58
rect 51 47 55 56
rect 51 45 53 47
rect 39 39 43 40
rect 39 37 40 39
rect 42 37 43 39
rect 7 29 8 31
rect 10 29 11 31
rect 7 24 11 29
rect 7 22 9 24
rect 11 22 19 24
rect 7 18 19 22
rect 39 31 43 37
rect 30 30 43 31
rect 30 28 35 30
rect 37 28 43 30
rect 30 26 43 28
rect 51 24 55 45
rect 66 63 79 64
rect 66 62 76 63
rect 66 60 70 62
rect 72 61 76 62
rect 78 61 79 63
rect 72 60 79 61
rect 66 58 79 60
rect 66 51 72 58
rect 95 47 99 56
rect 95 45 97 47
rect 83 39 87 40
rect 83 37 84 39
rect 86 37 87 39
rect 51 22 53 24
rect 55 22 63 24
rect 51 21 63 22
rect 51 19 56 21
rect 58 19 63 21
rect 51 18 63 19
rect 83 31 87 37
rect 74 30 87 31
rect 74 28 79 30
rect 81 28 87 30
rect 74 26 87 28
rect 95 24 99 45
rect 110 63 123 64
rect 110 62 120 63
rect 110 60 114 62
rect 116 61 120 62
rect 122 61 123 63
rect 116 60 123 61
rect 110 58 123 60
rect 110 51 116 58
rect 139 47 143 56
rect 139 45 141 47
rect 127 39 131 40
rect 127 37 128 39
rect 130 37 131 39
rect 95 22 97 24
rect 99 22 107 24
rect 95 21 107 22
rect 95 19 97 21
rect 99 19 107 21
rect 95 18 107 19
rect 127 31 131 37
rect 118 30 131 31
rect 118 28 123 30
rect 125 28 131 30
rect 118 26 131 28
rect 139 38 143 45
rect 154 63 167 64
rect 154 62 164 63
rect 154 60 158 62
rect 160 61 164 62
rect 166 61 167 63
rect 160 60 167 61
rect 154 58 167 60
rect 154 51 160 58
rect 183 47 187 56
rect 183 45 185 47
rect 139 36 140 38
rect 142 36 143 38
rect 139 24 143 36
rect 171 39 175 40
rect 171 37 172 39
rect 174 37 175 39
rect 139 22 141 24
rect 143 22 151 24
rect 139 18 151 22
rect 171 31 175 37
rect 162 30 175 31
rect 162 28 167 30
rect 169 28 175 30
rect 162 26 175 28
rect 183 29 187 45
rect 198 63 211 64
rect 198 62 208 63
rect 198 60 202 62
rect 204 61 208 62
rect 210 61 211 63
rect 204 60 211 61
rect 198 58 211 60
rect 198 51 204 58
rect 227 47 231 56
rect 227 45 229 47
rect 215 39 219 40
rect 215 37 216 39
rect 218 37 219 39
rect 183 27 184 29
rect 186 27 187 29
rect 183 24 187 27
rect 183 22 185 24
rect 187 22 195 24
rect 183 18 195 22
rect 215 31 219 37
rect 206 30 219 31
rect 206 28 211 30
rect 213 28 219 30
rect 206 26 219 28
rect 227 36 231 45
rect 242 63 255 64
rect 242 62 252 63
rect 242 60 246 62
rect 248 61 252 62
rect 254 61 255 63
rect 248 60 255 61
rect 242 58 255 60
rect 242 51 248 58
rect 271 47 275 56
rect 271 45 273 47
rect 227 34 228 36
rect 230 34 231 36
rect 259 39 263 40
rect 259 37 260 39
rect 262 37 263 39
rect 227 24 231 34
rect 227 22 229 24
rect 231 22 239 24
rect 227 18 239 22
rect 259 31 263 37
rect 250 30 263 31
rect 250 28 255 30
rect 257 28 263 30
rect 250 26 263 28
rect 271 24 275 45
rect 286 63 299 64
rect 286 62 296 63
rect 286 60 290 62
rect 292 61 296 62
rect 298 61 299 63
rect 292 60 299 61
rect 286 58 299 60
rect 286 51 292 58
rect 315 55 319 56
rect 315 53 316 55
rect 318 53 319 55
rect 315 47 319 53
rect 315 45 317 47
rect 303 39 307 40
rect 303 37 304 39
rect 306 37 307 39
rect 271 22 273 24
rect 275 22 283 24
rect 271 21 283 22
rect 271 19 272 21
rect 274 19 283 21
rect 271 18 283 19
rect 303 31 307 37
rect 294 30 307 31
rect 294 28 299 30
rect 301 28 307 30
rect 294 26 307 28
rect 315 24 319 45
rect 330 63 343 64
rect 330 62 340 63
rect 330 60 334 62
rect 336 61 340 62
rect 342 61 343 63
rect 336 60 343 61
rect 330 58 343 60
rect 330 51 336 58
rect 359 47 363 56
rect 359 45 361 47
rect 347 39 351 40
rect 347 37 348 39
rect 350 37 351 39
rect 315 22 317 24
rect 319 22 327 24
rect 315 18 327 22
rect 347 31 351 37
rect 338 30 351 31
rect 338 28 343 30
rect 345 28 351 30
rect 338 26 351 28
rect 359 24 363 45
rect 374 63 387 64
rect 374 62 384 63
rect 374 60 378 62
rect 380 61 384 62
rect 386 61 387 63
rect 380 60 387 61
rect 374 58 387 60
rect 374 51 380 58
rect 403 47 407 56
rect 403 45 405 47
rect 391 39 395 40
rect 391 37 392 39
rect 394 37 395 39
rect 359 22 361 24
rect 363 22 371 24
rect 359 21 371 22
rect 359 19 362 21
rect 364 19 371 21
rect 359 18 371 19
rect 391 31 395 37
rect 382 30 395 31
rect 382 28 387 30
rect 389 28 395 30
rect 382 26 395 28
rect 403 24 407 45
rect 418 63 431 64
rect 418 62 428 63
rect 418 60 422 62
rect 424 61 428 62
rect 430 61 431 63
rect 424 60 431 61
rect 418 58 431 60
rect 418 51 424 58
rect 447 47 451 56
rect 447 45 449 47
rect 435 39 439 40
rect 435 37 436 39
rect 438 37 439 39
rect 403 22 405 24
rect 407 22 415 24
rect 403 21 415 22
rect 403 19 405 21
rect 407 19 415 21
rect 403 18 415 19
rect 435 31 439 37
rect 426 30 439 31
rect 426 28 431 30
rect 433 28 439 30
rect 426 26 439 28
rect 447 30 451 45
rect 462 63 475 64
rect 462 62 472 63
rect 462 60 466 62
rect 468 61 472 62
rect 474 61 475 63
rect 468 60 475 61
rect 462 58 475 60
rect 462 51 468 58
rect 491 47 495 56
rect 491 45 493 47
rect 479 39 483 40
rect 479 37 480 39
rect 482 37 483 39
rect 447 28 448 30
rect 450 28 451 30
rect 447 24 451 28
rect 447 22 449 24
rect 451 22 459 24
rect 447 18 459 22
rect 479 31 483 37
rect 470 30 483 31
rect 470 28 475 30
rect 477 28 483 30
rect 470 26 483 28
rect 491 31 495 45
rect 506 63 519 64
rect 506 62 516 63
rect 506 60 510 62
rect 512 61 516 62
rect 518 61 519 63
rect 512 60 519 61
rect 506 58 519 60
rect 506 51 512 58
rect 535 47 539 56
rect 535 45 537 47
rect 523 39 527 40
rect 523 37 524 39
rect 526 37 527 39
rect 491 29 492 31
rect 494 29 495 31
rect 491 24 495 29
rect 491 22 493 24
rect 495 22 503 24
rect 491 18 503 22
rect 523 31 527 37
rect 514 30 527 31
rect 514 28 519 30
rect 521 28 527 30
rect 514 26 527 28
rect 535 30 539 45
rect 550 63 563 64
rect 550 62 560 63
rect 550 60 554 62
rect 556 61 560 62
rect 562 61 563 63
rect 556 60 563 61
rect 550 58 563 60
rect 550 51 556 58
rect 579 47 583 56
rect 579 45 581 47
rect 567 39 571 40
rect 567 37 568 39
rect 570 37 571 39
rect 535 28 536 30
rect 538 28 539 30
rect 535 24 539 28
rect 535 22 537 24
rect 539 22 547 24
rect 535 18 547 22
rect 567 31 571 37
rect 558 30 571 31
rect 558 28 563 30
rect 565 28 571 30
rect 558 26 571 28
rect 579 24 583 45
rect 594 63 607 64
rect 594 62 604 63
rect 594 60 598 62
rect 600 61 604 62
rect 606 61 607 63
rect 600 60 607 61
rect 594 58 607 60
rect 594 51 600 58
rect 623 47 627 56
rect 623 45 625 47
rect 611 39 615 40
rect 611 37 612 39
rect 614 37 615 39
rect 579 22 581 24
rect 583 22 591 24
rect 579 21 591 22
rect 579 19 580 21
rect 582 19 591 21
rect 579 18 591 19
rect 611 31 615 37
rect 602 30 615 31
rect 602 28 607 30
rect 609 28 615 30
rect 602 26 615 28
rect 623 24 627 45
rect 638 63 651 64
rect 638 62 648 63
rect 638 60 642 62
rect 644 61 648 62
rect 650 61 651 63
rect 644 60 651 61
rect 638 58 651 60
rect 638 51 644 58
rect 667 47 671 56
rect 667 45 669 47
rect 655 39 659 40
rect 655 37 656 39
rect 658 37 659 39
rect 623 22 625 24
rect 627 22 635 24
rect 623 21 635 22
rect 623 19 629 21
rect 631 19 635 21
rect 623 18 635 19
rect 655 31 659 37
rect 646 30 659 31
rect 646 28 651 30
rect 653 28 659 30
rect 646 26 659 28
rect 667 24 671 45
rect 682 63 695 64
rect 682 62 692 63
rect 682 60 686 62
rect 688 61 692 62
rect 694 61 695 63
rect 688 60 695 61
rect 682 58 695 60
rect 682 51 688 58
rect 699 39 703 40
rect 699 37 700 39
rect 702 37 703 39
rect 667 22 669 24
rect 671 22 679 24
rect 667 18 679 22
rect 699 31 703 37
rect 690 30 703 31
rect 690 28 695 30
rect 697 28 703 30
rect 690 26 703 28
rect -24 12 710 13
rect -24 10 10 12
rect 12 10 20 12
rect 22 10 54 12
rect 56 10 64 12
rect 66 10 98 12
rect 100 10 108 12
rect 110 10 142 12
rect 144 10 152 12
rect 154 10 186 12
rect 188 10 196 12
rect 198 10 230 12
rect 232 10 240 12
rect 242 10 274 12
rect 276 10 284 12
rect 286 10 318 12
rect 320 10 328 12
rect 330 10 362 12
rect 364 10 372 12
rect 374 10 406 12
rect 408 10 416 12
rect 418 10 450 12
rect 452 10 460 12
rect 462 10 494 12
rect 496 10 504 12
rect 506 10 538 12
rect 540 10 548 12
rect 550 10 582 12
rect 584 10 592 12
rect 594 10 626 12
rect 628 10 636 12
rect 638 10 670 12
rect 672 10 680 12
rect 682 10 710 12
rect -24 6 750 10
rect -24 4 -19 6
rect -17 5 745 6
rect -17 4 410 5
rect -24 0 410 4
rect -24 -2 195 0
rect 197 -2 223 0
rect 225 -2 410 0
rect -24 -3 410 -2
rect 479 -3 668 5
rect 707 4 745 5
rect 747 4 750 6
rect 707 0 750 4
rect 14 -10 36 -9
rect 14 -12 17 -10
rect 19 -12 36 -10
rect 14 -13 36 -12
rect 94 -10 99 -8
rect 94 -12 95 -10
rect 97 -12 99 -10
rect 14 -32 18 -13
rect 47 -17 51 -16
rect 47 -19 48 -17
rect 50 -19 51 -17
rect 14 -34 15 -32
rect 17 -33 18 -32
rect 17 -34 20 -33
rect 14 -35 20 -34
rect 14 -37 17 -35
rect 19 -37 20 -35
rect 14 -42 20 -37
rect 14 -44 17 -42
rect 19 -44 20 -42
rect 14 -46 20 -44
rect 47 -25 51 -19
rect 94 -14 99 -12
rect 63 -25 71 -24
rect 38 -26 53 -25
rect 38 -28 42 -26
rect 44 -28 49 -26
rect 51 -28 53 -26
rect 38 -29 53 -28
rect 63 -27 64 -25
rect 66 -26 71 -25
rect 66 -27 68 -26
rect 63 -28 68 -27
rect 70 -28 71 -26
rect 63 -30 71 -28
rect 63 -33 68 -30
rect 30 -37 68 -33
rect 95 -36 99 -14
rect 94 -38 99 -36
rect 94 -40 95 -38
rect 97 -40 99 -38
rect 94 -45 99 -40
rect 94 -47 95 -45
rect 97 -47 99 -45
rect 103 -10 125 -9
rect 103 -12 106 -10
rect 108 -12 125 -10
rect 103 -13 125 -12
rect 183 -10 188 -8
rect 183 -12 184 -10
rect 186 -12 188 -10
rect 103 -33 107 -13
rect 136 -17 140 -16
rect 136 -19 137 -17
rect 139 -19 140 -17
rect 103 -35 109 -33
rect 103 -37 106 -35
rect 108 -37 109 -35
rect 103 -39 109 -37
rect 103 -41 106 -39
rect 108 -41 109 -39
rect 103 -42 109 -41
rect 103 -44 106 -42
rect 108 -44 109 -42
rect 103 -46 109 -44
rect 136 -25 140 -19
rect 183 -14 188 -12
rect 184 -18 188 -14
rect 184 -20 185 -18
rect 187 -20 188 -18
rect 152 -25 160 -24
rect 127 -26 142 -25
rect 127 -28 131 -26
rect 133 -28 138 -26
rect 140 -28 142 -26
rect 127 -29 142 -28
rect 152 -27 153 -25
rect 155 -26 160 -25
rect 155 -27 157 -26
rect 152 -28 157 -27
rect 159 -28 160 -26
rect 152 -30 160 -28
rect 152 -33 157 -30
rect 119 -37 157 -33
rect 184 -36 188 -20
rect 223 -12 228 -8
rect 223 -14 224 -12
rect 226 -14 228 -12
rect 223 -16 228 -14
rect 183 -38 188 -36
rect 192 -25 196 -24
rect 192 -26 205 -25
rect 192 -28 197 -26
rect 199 -28 202 -26
rect 204 -28 205 -26
rect 192 -29 205 -28
rect 192 -38 196 -29
rect 200 -34 213 -33
rect 200 -36 207 -34
rect 209 -36 213 -34
rect 200 -37 213 -36
rect 200 -38 204 -37
rect 183 -40 184 -38
rect 186 -40 188 -38
rect 183 -45 188 -40
rect 94 -49 99 -47
rect 183 -47 184 -45
rect 186 -47 188 -45
rect 200 -40 201 -38
rect 203 -40 204 -38
rect 200 -46 204 -40
rect 224 -34 228 -16
rect 224 -36 225 -34
rect 227 -36 228 -34
rect 183 -49 188 -47
rect 224 -48 228 -36
rect 232 -10 254 -9
rect 232 -12 235 -10
rect 237 -12 254 -10
rect 232 -13 254 -12
rect 312 -10 317 -8
rect 312 -12 313 -10
rect 315 -12 317 -10
rect 232 -26 236 -13
rect 265 -18 269 -16
rect 265 -20 266 -18
rect 268 -20 269 -18
rect 232 -28 233 -26
rect 235 -28 236 -26
rect 232 -33 236 -28
rect 232 -35 238 -33
rect 232 -37 235 -35
rect 237 -37 238 -35
rect 232 -42 238 -37
rect 232 -44 235 -42
rect 237 -44 238 -42
rect 232 -46 238 -44
rect 265 -25 269 -20
rect 312 -14 317 -12
rect 256 -26 271 -25
rect 256 -28 260 -26
rect 262 -28 267 -26
rect 269 -28 271 -26
rect 256 -29 271 -28
rect 281 -26 289 -24
rect 281 -28 286 -26
rect 288 -28 289 -26
rect 281 -29 289 -28
rect 281 -31 282 -29
rect 284 -30 289 -29
rect 284 -31 286 -30
rect 281 -33 286 -31
rect 313 -24 317 -14
rect 313 -26 314 -24
rect 316 -26 317 -24
rect 248 -37 286 -33
rect 313 -36 317 -26
rect 312 -38 317 -36
rect 312 -40 313 -38
rect 315 -40 317 -38
rect 312 -45 317 -40
rect 86 -50 99 -49
rect 86 -52 89 -50
rect 91 -52 99 -50
rect 86 -53 99 -52
rect 175 -53 188 -49
rect 215 -50 224 -49
rect 226 -50 228 -48
rect 312 -47 313 -45
rect 315 -47 317 -45
rect 321 -10 343 -9
rect 321 -12 324 -10
rect 326 -12 343 -10
rect 321 -13 343 -12
rect 401 -10 406 -8
rect 401 -12 402 -10
rect 404 -12 406 -10
rect 321 -33 325 -13
rect 321 -35 327 -33
rect 321 -37 324 -35
rect 326 -37 327 -35
rect 321 -38 327 -37
rect 321 -40 322 -38
rect 324 -40 327 -38
rect 321 -42 327 -40
rect 321 -44 324 -42
rect 326 -44 327 -42
rect 321 -46 327 -44
rect 354 -25 358 -16
rect 401 -14 406 -12
rect 370 -25 378 -24
rect 345 -26 360 -25
rect 345 -28 346 -26
rect 348 -28 349 -26
rect 351 -28 356 -26
rect 358 -28 360 -26
rect 345 -29 360 -28
rect 370 -27 371 -25
rect 373 -26 378 -25
rect 373 -27 375 -26
rect 370 -28 375 -27
rect 377 -28 378 -26
rect 370 -30 378 -28
rect 370 -33 375 -30
rect 337 -37 375 -33
rect 402 -29 406 -14
rect 402 -31 403 -29
rect 405 -31 406 -29
rect 402 -36 406 -31
rect 401 -38 406 -36
rect 401 -40 402 -38
rect 404 -40 406 -38
rect 401 -45 406 -40
rect 312 -49 317 -47
rect 401 -47 402 -45
rect 404 -47 406 -45
rect 490 -10 512 -9
rect 490 -12 493 -10
rect 495 -12 512 -10
rect 490 -13 512 -12
rect 570 -10 575 -8
rect 570 -12 571 -10
rect 573 -12 575 -10
rect 490 -33 494 -13
rect 523 -17 527 -16
rect 523 -19 524 -17
rect 526 -19 527 -17
rect 490 -35 496 -33
rect 490 -37 493 -35
rect 495 -37 496 -35
rect 490 -39 496 -37
rect 490 -41 492 -39
rect 494 -41 496 -39
rect 490 -42 496 -41
rect 490 -44 493 -42
rect 495 -44 496 -42
rect 490 -46 496 -44
rect 523 -25 527 -19
rect 570 -14 575 -12
rect 514 -26 529 -25
rect 514 -28 518 -26
rect 520 -28 525 -26
rect 527 -28 529 -26
rect 514 -29 529 -28
rect 539 -26 547 -24
rect 539 -28 544 -26
rect 546 -28 547 -26
rect 539 -30 547 -28
rect 539 -33 544 -30
rect 506 -34 544 -33
rect 506 -36 536 -34
rect 538 -36 544 -34
rect 506 -37 544 -36
rect 571 -33 575 -14
rect 571 -35 572 -33
rect 574 -35 575 -33
rect 571 -36 575 -35
rect 570 -38 575 -36
rect 570 -40 571 -38
rect 573 -40 575 -38
rect 570 -45 575 -40
rect 401 -49 406 -47
rect 570 -47 571 -45
rect 573 -47 575 -45
rect 579 -10 601 -9
rect 579 -12 582 -10
rect 584 -12 601 -10
rect 579 -13 601 -12
rect 659 -10 664 -8
rect 659 -12 660 -10
rect 662 -12 664 -10
rect 579 -33 583 -13
rect 612 -17 616 -16
rect 612 -19 613 -17
rect 615 -19 616 -17
rect 579 -35 585 -33
rect 579 -37 582 -35
rect 584 -37 585 -35
rect 579 -39 585 -37
rect 579 -41 581 -39
rect 583 -41 585 -39
rect 579 -42 585 -41
rect 579 -44 582 -42
rect 584 -44 585 -42
rect 579 -46 585 -44
rect 612 -25 616 -19
rect 659 -14 664 -12
rect 628 -25 636 -24
rect 603 -26 618 -25
rect 603 -28 607 -26
rect 609 -28 614 -26
rect 616 -28 618 -26
rect 603 -29 618 -28
rect 628 -27 629 -25
rect 631 -26 636 -25
rect 631 -27 633 -26
rect 628 -28 633 -27
rect 635 -28 636 -26
rect 628 -30 636 -28
rect 628 -33 633 -30
rect 595 -37 633 -33
rect 660 -36 664 -14
rect 659 -38 664 -36
rect 659 -40 660 -38
rect 662 -40 664 -38
rect 659 -45 664 -40
rect 570 -49 575 -47
rect 659 -47 660 -45
rect 662 -47 664 -45
rect 659 -49 664 -47
rect 215 -53 228 -50
rect 304 -53 317 -49
rect 393 -53 406 -49
rect 562 -53 575 -49
rect 651 -53 664 -49
rect -1 -60 668 -59
rect -1 -62 223 -60
rect 225 -62 668 -60
rect -1 -63 739 -62
rect -21 -66 739 -63
rect -21 -68 -19 -66
rect -17 -68 732 -66
rect 734 -68 739 -66
rect -21 -71 739 -68
rect 3 -72 661 -71
rect 3 -74 188 -72
rect 190 -74 406 -72
rect 408 -74 624 -72
rect 626 -74 661 -72
rect 3 -75 661 -74
rect 7 -85 20 -81
rect 96 -85 109 -81
rect 185 -84 198 -81
rect 7 -87 12 -85
rect 7 -89 9 -87
rect 11 -89 12 -87
rect 96 -87 101 -85
rect 7 -94 12 -89
rect 7 -96 9 -94
rect 11 -96 12 -94
rect 7 -98 12 -96
rect 7 -103 11 -98
rect 7 -105 8 -103
rect 10 -105 11 -103
rect 7 -120 11 -105
rect 38 -98 76 -97
rect 38 -100 56 -98
rect 58 -100 76 -98
rect 38 -101 76 -100
rect 38 -104 43 -101
rect 35 -106 43 -104
rect 35 -108 36 -106
rect 38 -108 43 -106
rect 35 -110 43 -108
rect 53 -106 68 -105
rect 53 -108 55 -106
rect 57 -108 62 -106
rect 64 -108 68 -106
rect 53 -109 68 -108
rect 55 -111 59 -109
rect 86 -90 92 -88
rect 86 -92 87 -90
rect 89 -92 92 -90
rect 86 -94 92 -92
rect 86 -96 89 -94
rect 91 -96 92 -94
rect 86 -97 92 -96
rect 86 -99 87 -97
rect 89 -99 92 -97
rect 86 -101 92 -99
rect 55 -113 56 -111
rect 58 -113 59 -111
rect 7 -122 12 -120
rect 55 -118 59 -113
rect 88 -121 92 -101
rect 7 -124 9 -122
rect 11 -124 12 -122
rect 7 -126 12 -124
rect 70 -122 92 -121
rect 70 -124 87 -122
rect 89 -124 92 -122
rect 70 -125 92 -124
rect 96 -89 98 -87
rect 100 -89 101 -87
rect 185 -86 187 -84
rect 189 -85 198 -84
rect 225 -85 238 -81
rect 314 -85 327 -81
rect 403 -84 416 -81
rect 96 -94 101 -89
rect 96 -96 98 -94
rect 100 -96 101 -94
rect 96 -98 101 -96
rect 96 -119 100 -98
rect 127 -101 165 -97
rect 127 -103 132 -101
rect 127 -104 129 -103
rect 124 -105 129 -104
rect 131 -105 132 -103
rect 124 -106 132 -105
rect 124 -108 125 -106
rect 127 -108 132 -106
rect 124 -110 132 -108
rect 142 -106 157 -105
rect 142 -108 144 -106
rect 146 -108 151 -106
rect 153 -108 157 -106
rect 142 -109 157 -108
rect 144 -111 148 -109
rect 175 -90 181 -88
rect 175 -92 176 -90
rect 178 -92 181 -90
rect 175 -97 181 -92
rect 175 -99 176 -97
rect 178 -99 181 -97
rect 175 -101 181 -99
rect 177 -106 181 -101
rect 177 -108 178 -106
rect 180 -108 181 -106
rect 144 -113 145 -111
rect 147 -113 148 -111
rect 96 -121 97 -119
rect 99 -120 100 -119
rect 99 -121 101 -120
rect 96 -122 101 -121
rect 144 -118 148 -113
rect 177 -121 181 -108
rect 96 -124 98 -122
rect 100 -124 101 -122
rect 96 -126 101 -124
rect 159 -122 181 -121
rect 159 -124 176 -122
rect 178 -124 181 -122
rect 159 -125 181 -124
rect 185 -114 189 -86
rect 225 -87 230 -85
rect 185 -116 186 -114
rect 188 -116 189 -114
rect 209 -94 213 -88
rect 209 -96 210 -94
rect 212 -96 213 -94
rect 225 -89 227 -87
rect 229 -89 230 -87
rect 314 -87 319 -85
rect 225 -94 230 -89
rect 225 -96 227 -94
rect 229 -96 230 -94
rect 209 -97 213 -96
rect 200 -98 213 -97
rect 200 -100 204 -98
rect 206 -100 213 -98
rect 200 -101 213 -100
rect 217 -105 221 -96
rect 208 -106 221 -105
rect 208 -108 209 -106
rect 211 -108 214 -106
rect 216 -108 221 -106
rect 208 -109 221 -108
rect 217 -110 221 -109
rect 225 -98 230 -96
rect 225 -103 229 -98
rect 225 -105 226 -103
rect 228 -105 229 -103
rect 185 -118 189 -116
rect 185 -120 190 -118
rect 185 -122 187 -120
rect 189 -122 190 -120
rect 185 -126 190 -122
rect 225 -120 229 -105
rect 256 -98 294 -97
rect 256 -100 258 -98
rect 260 -100 294 -98
rect 256 -101 294 -100
rect 256 -104 261 -101
rect 253 -106 261 -104
rect 253 -108 254 -106
rect 256 -108 261 -106
rect 253 -110 261 -108
rect 271 -106 286 -105
rect 271 -108 273 -106
rect 275 -108 280 -106
rect 282 -108 286 -106
rect 271 -109 286 -108
rect 273 -111 277 -109
rect 304 -90 310 -88
rect 304 -92 305 -90
rect 307 -92 310 -90
rect 304 -94 310 -92
rect 304 -96 307 -94
rect 309 -96 310 -94
rect 304 -97 310 -96
rect 304 -99 305 -97
rect 307 -99 310 -97
rect 304 -101 310 -99
rect 273 -113 274 -111
rect 276 -113 277 -111
rect 225 -122 230 -120
rect 273 -118 277 -113
rect 306 -121 310 -101
rect 225 -124 227 -122
rect 229 -124 230 -122
rect 225 -126 230 -124
rect 288 -122 310 -121
rect 288 -124 305 -122
rect 307 -124 310 -122
rect 288 -125 310 -124
rect 314 -89 316 -87
rect 318 -89 319 -87
rect 403 -86 405 -84
rect 407 -85 416 -84
rect 443 -85 456 -81
rect 532 -85 545 -81
rect 621 -84 634 -81
rect 314 -94 319 -89
rect 314 -96 316 -94
rect 318 -96 319 -94
rect 314 -98 319 -96
rect 314 -117 318 -98
rect 345 -101 383 -97
rect 345 -103 350 -101
rect 345 -104 347 -103
rect 342 -105 347 -104
rect 349 -105 350 -103
rect 342 -106 350 -105
rect 342 -108 343 -106
rect 345 -108 350 -106
rect 342 -110 350 -108
rect 360 -106 375 -105
rect 360 -108 362 -106
rect 364 -108 369 -106
rect 371 -108 375 -106
rect 360 -109 375 -108
rect 362 -111 366 -109
rect 393 -90 399 -88
rect 393 -92 394 -90
rect 396 -92 399 -90
rect 393 -97 399 -92
rect 393 -99 394 -97
rect 396 -99 399 -97
rect 393 -101 399 -99
rect 395 -106 399 -101
rect 395 -108 396 -106
rect 398 -108 399 -106
rect 362 -113 363 -111
rect 365 -113 366 -111
rect 314 -119 315 -117
rect 317 -119 318 -117
rect 314 -120 318 -119
rect 314 -122 319 -120
rect 362 -118 366 -113
rect 395 -121 399 -108
rect 314 -124 316 -122
rect 318 -124 319 -122
rect 314 -126 319 -124
rect 377 -122 399 -121
rect 377 -124 394 -122
rect 396 -124 399 -122
rect 377 -125 399 -124
rect 403 -112 407 -86
rect 443 -87 448 -85
rect 403 -114 404 -112
rect 406 -114 407 -112
rect 403 -118 407 -114
rect 427 -94 431 -88
rect 427 -96 428 -94
rect 430 -96 431 -94
rect 443 -89 445 -87
rect 447 -89 448 -87
rect 532 -87 537 -85
rect 443 -94 448 -89
rect 443 -96 445 -94
rect 447 -96 448 -94
rect 427 -97 431 -96
rect 418 -98 431 -97
rect 418 -100 422 -98
rect 424 -100 431 -98
rect 418 -101 431 -100
rect 435 -105 439 -96
rect 426 -106 439 -105
rect 426 -108 427 -106
rect 429 -108 432 -106
rect 434 -108 439 -106
rect 426 -109 439 -108
rect 435 -110 439 -109
rect 443 -98 448 -96
rect 443 -103 447 -98
rect 443 -105 444 -103
rect 446 -105 447 -103
rect 403 -120 408 -118
rect 403 -122 405 -120
rect 407 -122 408 -120
rect 403 -126 408 -122
rect 443 -120 447 -105
rect 474 -98 512 -97
rect 474 -100 484 -98
rect 486 -100 512 -98
rect 474 -101 512 -100
rect 474 -104 479 -101
rect 471 -106 479 -104
rect 471 -108 472 -106
rect 474 -108 479 -106
rect 471 -110 479 -108
rect 489 -106 504 -105
rect 489 -108 491 -106
rect 493 -108 498 -106
rect 500 -108 504 -106
rect 489 -109 504 -108
rect 491 -111 495 -109
rect 522 -90 528 -88
rect 522 -92 523 -90
rect 525 -92 528 -90
rect 522 -94 528 -92
rect 522 -96 525 -94
rect 527 -96 528 -94
rect 522 -97 528 -96
rect 522 -99 523 -97
rect 525 -99 528 -97
rect 522 -101 528 -99
rect 491 -113 492 -111
rect 494 -113 495 -111
rect 443 -122 448 -120
rect 491 -118 495 -113
rect 524 -121 528 -101
rect 443 -124 445 -122
rect 447 -124 448 -122
rect 443 -126 448 -124
rect 506 -122 528 -121
rect 506 -124 523 -122
rect 525 -124 528 -122
rect 506 -125 528 -124
rect 532 -89 534 -87
rect 536 -89 537 -87
rect 621 -86 623 -84
rect 625 -85 634 -84
rect 532 -94 537 -89
rect 532 -96 534 -94
rect 536 -96 537 -94
rect 532 -98 537 -96
rect 532 -120 536 -98
rect 563 -101 601 -97
rect 563 -103 568 -101
rect 563 -104 565 -103
rect 560 -105 565 -104
rect 567 -105 568 -103
rect 560 -106 568 -105
rect 560 -108 561 -106
rect 563 -108 568 -106
rect 560 -110 568 -108
rect 578 -106 593 -105
rect 578 -108 580 -106
rect 582 -108 587 -106
rect 589 -108 593 -106
rect 578 -109 593 -108
rect 580 -111 584 -109
rect 611 -90 617 -88
rect 611 -92 612 -90
rect 614 -92 617 -90
rect 611 -97 617 -92
rect 611 -99 612 -97
rect 614 -99 617 -97
rect 611 -101 617 -99
rect 613 -106 617 -101
rect 613 -108 614 -106
rect 616 -108 617 -106
rect 580 -113 581 -111
rect 583 -113 584 -111
rect 532 -122 537 -120
rect 580 -118 584 -113
rect 613 -121 617 -108
rect 532 -124 534 -122
rect 536 -124 537 -122
rect 532 -126 537 -124
rect 595 -122 617 -121
rect 595 -124 612 -122
rect 614 -124 617 -122
rect 595 -125 617 -124
rect 621 -115 625 -86
rect 621 -117 622 -115
rect 624 -117 625 -115
rect 645 -94 649 -88
rect 645 -96 646 -94
rect 648 -96 649 -94
rect 645 -97 649 -96
rect 636 -98 649 -97
rect 636 -100 640 -98
rect 642 -100 649 -98
rect 636 -101 649 -100
rect 653 -105 657 -96
rect 644 -106 657 -105
rect 644 -108 645 -106
rect 647 -108 650 -106
rect 652 -108 657 -106
rect 644 -109 657 -108
rect 653 -110 657 -109
rect 621 -118 625 -117
rect 621 -120 626 -118
rect 621 -122 623 -120
rect 625 -122 626 -120
rect 621 -126 626 -122
rect -30 -132 719 -131
rect -30 -134 188 -132
rect 190 -134 216 -132
rect 218 -134 406 -132
rect 408 -134 434 -132
rect 436 -134 624 -132
rect 626 -134 652 -132
rect 654 -134 719 -132
rect -30 -136 -28 -134
rect -26 -136 755 -134
rect -30 -138 755 -136
rect -30 -139 750 -138
rect 228 -140 750 -139
rect 752 -140 755 -138
rect 228 -144 755 -140
rect 228 -146 235 -144
rect 237 -146 263 -144
rect 265 -146 479 -144
rect 481 -146 507 -144
rect 509 -146 716 -144
rect 228 -147 716 -146
rect 263 -156 268 -152
rect 263 -158 264 -156
rect 266 -158 268 -156
rect 263 -160 268 -158
rect 232 -169 236 -168
rect 232 -170 245 -169
rect 232 -172 237 -170
rect 239 -172 242 -170
rect 244 -172 245 -170
rect 232 -173 245 -172
rect 232 -182 236 -173
rect 240 -178 253 -177
rect 240 -180 247 -178
rect 249 -180 253 -178
rect 240 -181 253 -180
rect 240 -182 244 -181
rect 240 -184 241 -182
rect 243 -184 244 -182
rect 240 -190 244 -184
rect 264 -177 268 -160
rect 264 -179 265 -177
rect 267 -179 268 -177
rect 264 -192 268 -179
rect 283 -154 305 -153
rect 283 -156 286 -154
rect 288 -156 305 -154
rect 283 -157 305 -156
rect 363 -154 368 -152
rect 363 -156 364 -154
rect 366 -156 368 -154
rect 283 -170 287 -157
rect 316 -161 320 -160
rect 316 -163 317 -161
rect 319 -163 320 -161
rect 283 -172 284 -170
rect 286 -172 287 -170
rect 283 -177 287 -172
rect 283 -179 289 -177
rect 283 -181 286 -179
rect 288 -181 289 -179
rect 283 -186 289 -181
rect 283 -188 286 -186
rect 288 -188 289 -186
rect 283 -190 289 -188
rect 316 -169 320 -163
rect 363 -158 368 -156
rect 307 -170 322 -169
rect 307 -172 311 -170
rect 313 -172 318 -170
rect 320 -172 322 -170
rect 307 -173 322 -172
rect 332 -170 340 -168
rect 332 -172 337 -170
rect 339 -172 340 -170
rect 332 -173 340 -172
rect 332 -175 333 -173
rect 335 -174 340 -173
rect 335 -175 337 -174
rect 332 -177 337 -175
rect 299 -181 337 -177
rect 364 -180 368 -158
rect 363 -182 368 -180
rect 363 -184 364 -182
rect 366 -184 368 -182
rect 363 -189 368 -184
rect 255 -194 264 -193
rect 266 -194 268 -192
rect 363 -191 364 -189
rect 366 -191 368 -189
rect 383 -154 405 -153
rect 383 -156 386 -154
rect 388 -156 405 -154
rect 383 -157 405 -156
rect 463 -154 468 -152
rect 463 -156 464 -154
rect 466 -156 468 -154
rect 383 -177 387 -157
rect 416 -161 420 -160
rect 416 -163 417 -161
rect 419 -163 420 -161
rect 383 -179 389 -177
rect 383 -181 386 -179
rect 388 -181 389 -179
rect 383 -182 389 -181
rect 383 -184 384 -182
rect 386 -184 389 -182
rect 383 -186 389 -184
rect 383 -188 386 -186
rect 388 -188 389 -186
rect 383 -190 389 -188
rect 416 -169 420 -163
rect 463 -158 468 -156
rect 407 -170 422 -169
rect 407 -172 411 -170
rect 413 -172 418 -170
rect 420 -172 422 -170
rect 407 -173 422 -172
rect 432 -170 440 -168
rect 432 -172 437 -170
rect 439 -172 440 -170
rect 432 -174 440 -172
rect 432 -177 437 -174
rect 399 -178 437 -177
rect 399 -180 434 -178
rect 436 -180 437 -178
rect 399 -181 437 -180
rect 464 -173 468 -158
rect 507 -156 512 -152
rect 507 -158 508 -156
rect 510 -158 512 -156
rect 507 -160 512 -158
rect 464 -175 465 -173
rect 467 -175 468 -173
rect 464 -180 468 -175
rect 463 -182 468 -180
rect 476 -169 480 -168
rect 476 -170 489 -169
rect 476 -172 481 -170
rect 483 -172 486 -170
rect 488 -172 489 -170
rect 476 -173 489 -172
rect 476 -182 480 -173
rect 484 -178 497 -177
rect 484 -180 491 -178
rect 493 -180 497 -178
rect 484 -181 497 -180
rect 484 -182 488 -181
rect 463 -184 464 -182
rect 466 -184 468 -182
rect 463 -189 468 -184
rect 363 -193 368 -191
rect 463 -191 464 -189
rect 466 -191 468 -189
rect 484 -184 485 -182
rect 487 -184 488 -182
rect 484 -190 488 -184
rect 463 -193 468 -191
rect 508 -192 512 -160
rect 527 -154 549 -153
rect 527 -156 530 -154
rect 532 -156 549 -154
rect 527 -157 549 -156
rect 607 -154 612 -152
rect 607 -156 608 -154
rect 610 -156 612 -154
rect 527 -170 531 -157
rect 560 -162 564 -160
rect 560 -164 561 -162
rect 563 -164 564 -162
rect 527 -172 528 -170
rect 530 -172 531 -170
rect 527 -177 531 -172
rect 527 -179 533 -177
rect 527 -181 530 -179
rect 532 -181 533 -179
rect 527 -186 533 -181
rect 527 -188 530 -186
rect 532 -188 533 -186
rect 527 -190 533 -188
rect 560 -169 564 -164
rect 607 -158 612 -156
rect 551 -170 566 -169
rect 551 -172 555 -170
rect 557 -172 562 -170
rect 564 -172 566 -170
rect 551 -173 566 -172
rect 576 -170 584 -168
rect 576 -172 581 -170
rect 583 -172 584 -170
rect 576 -173 584 -172
rect 576 -175 577 -173
rect 579 -174 584 -173
rect 579 -175 581 -174
rect 576 -177 581 -175
rect 543 -181 581 -177
rect 608 -180 612 -158
rect 607 -182 612 -180
rect 607 -184 608 -182
rect 610 -184 612 -182
rect 607 -189 612 -184
rect 255 -197 268 -194
rect 355 -197 368 -193
rect 455 -197 468 -193
rect 499 -194 508 -193
rect 510 -194 512 -192
rect 607 -191 608 -189
rect 610 -191 612 -189
rect 627 -154 649 -153
rect 627 -156 630 -154
rect 632 -156 649 -154
rect 627 -157 649 -156
rect 707 -154 712 -152
rect 707 -156 708 -154
rect 710 -156 712 -154
rect 627 -177 631 -157
rect 660 -161 664 -160
rect 660 -163 661 -161
rect 663 -163 664 -161
rect 627 -179 633 -177
rect 627 -181 630 -179
rect 632 -181 633 -179
rect 627 -182 633 -181
rect 627 -184 628 -182
rect 630 -184 633 -182
rect 627 -186 633 -184
rect 627 -188 630 -186
rect 632 -188 633 -186
rect 627 -190 633 -188
rect 660 -169 664 -163
rect 707 -158 712 -156
rect 651 -170 666 -169
rect 651 -172 655 -170
rect 657 -172 662 -170
rect 664 -172 666 -170
rect 651 -173 666 -172
rect 676 -170 684 -168
rect 676 -172 681 -170
rect 683 -172 684 -170
rect 676 -174 684 -172
rect 676 -177 681 -174
rect 643 -178 681 -177
rect 643 -180 669 -178
rect 671 -180 681 -178
rect 643 -181 681 -180
rect 708 -173 712 -158
rect 708 -175 709 -173
rect 711 -175 712 -173
rect 708 -180 712 -175
rect 707 -182 712 -180
rect 707 -184 708 -182
rect 710 -184 712 -182
rect 707 -189 712 -184
rect 607 -193 612 -191
rect 707 -191 708 -189
rect 710 -191 712 -189
rect 707 -193 712 -191
rect 499 -196 500 -194
rect 502 -196 512 -194
rect 499 -197 512 -196
rect 599 -197 612 -193
rect 699 -197 712 -193
rect -1 -204 742 -203
rect -1 -206 263 -204
rect 265 -206 507 -204
rect 509 -206 742 -204
rect -1 -207 737 -206
rect -22 -208 737 -207
rect 739 -208 742 -206
rect -22 -210 742 -208
rect -22 -212 -20 -210
rect -18 -211 742 -210
rect -18 -212 488 -211
rect -22 -215 488 -212
rect 3 -216 488 -215
rect 3 -218 210 -216
rect 212 -218 451 -216
rect 453 -218 488 -216
rect 3 -219 488 -218
rect 7 -229 20 -225
rect 107 -229 120 -225
rect 207 -228 220 -225
rect 7 -231 12 -229
rect 7 -233 9 -231
rect 11 -233 12 -231
rect 107 -231 112 -229
rect 7 -238 12 -233
rect 7 -240 9 -238
rect 11 -240 12 -238
rect 7 -242 12 -240
rect 7 -247 11 -242
rect 7 -249 8 -247
rect 10 -249 11 -247
rect 7 -264 11 -249
rect 38 -242 76 -241
rect 38 -244 67 -242
rect 69 -244 76 -242
rect 38 -245 76 -244
rect 38 -248 43 -245
rect 35 -250 43 -248
rect 35 -252 36 -250
rect 38 -252 43 -250
rect 35 -254 43 -252
rect 53 -250 68 -249
rect 53 -252 55 -250
rect 57 -252 62 -250
rect 64 -252 68 -250
rect 53 -253 68 -252
rect 55 -255 59 -253
rect 86 -234 92 -232
rect 86 -236 87 -234
rect 89 -236 92 -234
rect 86 -238 92 -236
rect 86 -240 89 -238
rect 91 -240 92 -238
rect 86 -241 92 -240
rect 86 -243 87 -241
rect 89 -243 92 -241
rect 86 -245 92 -243
rect 55 -257 56 -255
rect 58 -257 59 -255
rect 7 -266 12 -264
rect 55 -262 59 -257
rect 88 -265 92 -245
rect 7 -268 9 -266
rect 11 -268 12 -266
rect 7 -270 12 -268
rect 70 -266 92 -265
rect 70 -268 87 -266
rect 89 -268 92 -266
rect 70 -269 92 -268
rect 107 -233 109 -231
rect 111 -233 112 -231
rect 207 -230 209 -228
rect 211 -229 220 -228
rect 248 -229 261 -225
rect 348 -229 361 -225
rect 448 -228 461 -225
rect 107 -238 112 -233
rect 107 -240 109 -238
rect 111 -240 112 -238
rect 107 -242 112 -240
rect 107 -264 111 -242
rect 138 -245 176 -241
rect 138 -247 143 -245
rect 138 -248 140 -247
rect 135 -249 140 -248
rect 142 -249 143 -247
rect 135 -250 143 -249
rect 135 -252 136 -250
rect 138 -252 143 -250
rect 135 -254 143 -252
rect 153 -250 168 -249
rect 153 -252 155 -250
rect 157 -252 162 -250
rect 164 -252 168 -250
rect 153 -253 168 -252
rect 155 -255 159 -253
rect 186 -234 192 -232
rect 186 -236 187 -234
rect 189 -236 192 -234
rect 186 -241 192 -236
rect 186 -243 187 -241
rect 189 -243 192 -241
rect 186 -245 192 -243
rect 188 -250 192 -245
rect 188 -252 189 -250
rect 191 -252 192 -250
rect 155 -257 156 -255
rect 158 -257 159 -255
rect 107 -266 112 -264
rect 155 -262 159 -257
rect 188 -265 192 -252
rect 107 -268 109 -266
rect 111 -268 112 -266
rect 107 -270 112 -268
rect 170 -266 192 -265
rect 170 -268 187 -266
rect 189 -268 192 -266
rect 170 -269 192 -268
rect 207 -258 211 -230
rect 248 -231 253 -229
rect 207 -260 208 -258
rect 210 -260 211 -258
rect 231 -238 235 -232
rect 231 -240 232 -238
rect 234 -240 235 -238
rect 248 -233 250 -231
rect 252 -233 253 -231
rect 348 -231 353 -229
rect 248 -238 253 -233
rect 248 -240 250 -238
rect 252 -240 253 -238
rect 231 -241 235 -240
rect 222 -242 235 -241
rect 222 -244 226 -242
rect 228 -244 235 -242
rect 222 -245 235 -244
rect 239 -249 243 -240
rect 230 -250 243 -249
rect 230 -252 231 -250
rect 233 -252 236 -250
rect 238 -252 243 -250
rect 230 -253 243 -252
rect 239 -254 243 -253
rect 248 -242 253 -240
rect 248 -247 252 -242
rect 248 -249 249 -247
rect 251 -249 252 -247
rect 207 -262 211 -260
rect 207 -264 212 -262
rect 207 -266 209 -264
rect 211 -266 212 -264
rect 207 -270 212 -266
rect 248 -264 252 -249
rect 279 -242 317 -241
rect 279 -244 280 -242
rect 282 -244 317 -242
rect 279 -245 317 -244
rect 279 -248 284 -245
rect 276 -250 284 -248
rect 276 -252 277 -250
rect 279 -252 284 -250
rect 276 -254 284 -252
rect 294 -250 309 -249
rect 294 -252 296 -250
rect 298 -252 303 -250
rect 305 -252 309 -250
rect 294 -253 309 -252
rect 248 -266 253 -264
rect 296 -258 300 -253
rect 327 -234 333 -232
rect 327 -236 328 -234
rect 330 -236 333 -234
rect 327 -238 333 -236
rect 327 -240 330 -238
rect 332 -240 333 -238
rect 327 -241 333 -240
rect 327 -243 328 -241
rect 330 -243 333 -241
rect 327 -245 333 -243
rect 296 -260 297 -258
rect 299 -260 300 -258
rect 296 -262 300 -260
rect 329 -265 333 -245
rect 248 -268 250 -266
rect 252 -268 253 -266
rect 248 -270 253 -268
rect 311 -266 333 -265
rect 311 -268 328 -266
rect 330 -268 333 -266
rect 311 -269 333 -268
rect 348 -233 350 -231
rect 352 -233 353 -231
rect 448 -230 450 -228
rect 452 -229 461 -228
rect 348 -238 353 -233
rect 348 -240 350 -238
rect 352 -240 353 -238
rect 348 -242 353 -240
rect 348 -264 352 -242
rect 379 -245 417 -241
rect 379 -247 384 -245
rect 379 -248 381 -247
rect 376 -249 381 -248
rect 383 -249 384 -247
rect 376 -250 384 -249
rect 376 -252 377 -250
rect 379 -252 384 -250
rect 376 -254 384 -252
rect 394 -250 409 -249
rect 394 -252 396 -250
rect 398 -252 403 -250
rect 405 -252 409 -250
rect 394 -253 409 -252
rect 348 -266 353 -264
rect 396 -259 400 -253
rect 427 -234 433 -232
rect 427 -236 428 -234
rect 430 -236 433 -234
rect 427 -241 433 -236
rect 427 -243 428 -241
rect 430 -243 433 -241
rect 427 -245 433 -243
rect 429 -250 433 -245
rect 429 -252 430 -250
rect 432 -252 433 -250
rect 396 -261 397 -259
rect 399 -261 400 -259
rect 396 -262 400 -261
rect 429 -265 433 -252
rect 348 -268 350 -266
rect 352 -268 353 -266
rect 348 -270 353 -268
rect 411 -266 433 -265
rect 411 -268 428 -266
rect 430 -268 433 -266
rect 411 -269 433 -268
rect 448 -262 452 -230
rect 472 -238 476 -232
rect 472 -240 473 -238
rect 475 -240 476 -238
rect 472 -241 476 -240
rect 463 -242 476 -241
rect 463 -244 467 -242
rect 469 -244 476 -242
rect 463 -245 476 -244
rect 480 -249 484 -240
rect 471 -250 484 -249
rect 471 -252 472 -250
rect 474 -252 477 -250
rect 479 -252 484 -250
rect 471 -253 484 -252
rect 480 -254 484 -253
rect 448 -264 453 -262
rect 448 -266 450 -264
rect 452 -266 453 -264
rect 448 -270 453 -266
rect -33 -276 726 -275
rect -33 -278 210 -276
rect 212 -278 238 -276
rect 240 -278 451 -276
rect 453 -278 479 -276
rect 481 -278 726 -276
rect -33 -280 -31 -278
rect -29 -280 719 -278
rect 721 -280 726 -278
rect -33 -282 726 -280
rect 3 -283 726 -282
<< alu2 >>
rect 39 142 43 143
rect 39 140 40 142
rect 42 140 43 142
rect 31 134 35 135
rect 31 132 32 134
rect 34 132 35 134
rect -22 74 -15 77
rect -22 72 -19 74
rect -17 72 -15 74
rect -22 69 -15 72
rect 31 63 35 132
rect 31 61 32 63
rect 34 61 35 63
rect 31 60 35 61
rect 39 39 43 140
rect 83 142 87 143
rect 83 140 84 142
rect 86 140 87 142
rect 75 118 79 119
rect 75 116 76 118
rect 78 116 79 118
rect 75 63 79 116
rect 75 61 76 63
rect 78 61 79 63
rect 75 60 79 61
rect 83 39 87 140
rect 171 142 175 143
rect 171 140 172 142
rect 174 140 175 142
rect 119 134 123 135
rect 119 132 120 134
rect 122 132 123 134
rect 119 63 123 132
rect 119 61 120 63
rect 122 61 123 63
rect 119 60 123 61
rect 127 126 131 127
rect 127 124 128 126
rect 130 124 131 126
rect 39 37 40 39
rect 42 37 43 39
rect 39 36 43 37
rect 47 38 51 39
rect 47 36 48 38
rect 50 36 51 38
rect 83 37 84 39
rect 86 37 87 39
rect 83 36 87 37
rect 127 39 131 124
rect 163 102 167 103
rect 163 100 164 102
rect 166 100 167 102
rect 163 63 167 100
rect 163 61 164 63
rect 166 61 167 63
rect 163 60 167 61
rect 152 55 156 56
rect 152 53 153 55
rect 155 53 156 55
rect 127 37 128 39
rect 130 37 131 39
rect 127 36 131 37
rect 139 38 143 39
rect 139 36 140 38
rect 142 36 143 38
rect -1 31 3 32
rect -1 29 0 31
rect 2 29 3 31
rect -24 6 -12 13
rect -24 4 -19 6
rect -17 4 -12 6
rect -24 -3 -12 4
rect -21 -66 -15 -63
rect -21 -68 -19 -66
rect -17 -68 -15 -66
rect -21 -71 -15 -68
rect -30 -134 -24 -131
rect -30 -136 -28 -134
rect -26 -136 -24 -134
rect -30 -139 -24 -136
rect -22 -210 -15 -207
rect -22 -212 -20 -210
rect -18 -212 -15 -210
rect -22 -215 -15 -212
rect -33 -278 -27 -275
rect -33 -280 -31 -278
rect -29 -280 -27 -278
rect -33 -282 -27 -280
rect -1 -280 3 29
rect 7 31 11 32
rect 7 29 8 31
rect 10 29 11 31
rect 7 28 11 29
rect 47 -17 51 36
rect 139 35 143 36
rect 63 29 67 30
rect 63 27 64 29
rect 66 27 67 29
rect 47 -19 48 -17
rect 50 -19 51 -17
rect 47 -20 51 -19
rect 55 21 59 22
rect 55 19 56 21
rect 58 19 59 21
rect 14 -32 19 -31
rect 14 -34 15 -32
rect 17 -34 19 -32
rect 14 -35 19 -34
rect 55 -98 59 19
rect 63 -25 67 27
rect 96 21 100 22
rect 96 19 97 21
rect 99 19 100 21
rect 63 -27 64 -25
rect 66 -27 67 -25
rect 63 -29 67 -27
rect 88 -5 92 -4
rect 88 -7 89 -5
rect 91 -7 92 -5
rect 88 -50 92 -7
rect 88 -52 89 -50
rect 91 -52 92 -50
rect 88 -53 92 -52
rect 88 -94 92 -93
rect 88 -96 89 -94
rect 91 -96 92 -94
rect 88 -97 92 -96
rect 55 -100 56 -98
rect 58 -100 59 -98
rect 55 -101 59 -100
rect 7 -103 11 -102
rect 7 -105 8 -103
rect 10 -105 11 -103
rect 7 -106 11 -105
rect 55 -111 59 -110
rect 55 -113 56 -111
rect 58 -113 59 -111
rect 55 -114 59 -113
rect 96 -111 100 19
rect 136 21 140 22
rect 136 19 137 21
rect 139 19 140 21
rect 136 -17 140 19
rect 136 -19 137 -17
rect 139 -19 140 -17
rect 136 -20 140 -19
rect 152 -25 156 53
rect 171 39 175 140
rect 303 142 307 143
rect 303 140 304 142
rect 306 140 307 142
rect 251 134 255 135
rect 251 132 252 134
rect 254 132 255 134
rect 215 126 219 127
rect 215 124 216 126
rect 218 124 219 126
rect 207 118 211 119
rect 207 116 208 118
rect 210 116 211 118
rect 207 63 211 116
rect 207 61 208 63
rect 210 61 211 63
rect 207 60 211 61
rect 171 37 172 39
rect 174 37 175 39
rect 171 36 175 37
rect 215 39 219 124
rect 251 63 255 132
rect 251 61 252 63
rect 254 61 255 63
rect 251 60 255 61
rect 259 110 263 111
rect 259 108 260 110
rect 262 108 263 110
rect 215 37 216 39
rect 218 37 219 39
rect 259 39 263 108
rect 295 86 299 87
rect 295 84 296 86
rect 298 84 299 86
rect 295 63 299 84
rect 295 61 296 63
rect 298 61 299 63
rect 295 60 299 61
rect 259 37 260 39
rect 262 37 263 39
rect 215 36 219 37
rect 227 36 231 37
rect 259 36 263 37
rect 303 39 307 140
rect 427 134 431 135
rect 427 132 428 134
rect 430 132 431 134
rect 347 126 351 127
rect 347 124 348 126
rect 350 124 351 126
rect 339 102 343 103
rect 339 100 340 102
rect 342 100 343 102
rect 339 63 343 100
rect 339 61 340 63
rect 342 61 343 63
rect 339 60 343 61
rect 315 55 319 56
rect 315 53 316 55
rect 318 53 319 55
rect 315 52 319 53
rect 303 37 304 39
rect 306 37 307 39
rect 303 36 307 37
rect 347 39 351 124
rect 383 118 387 119
rect 383 116 384 118
rect 386 116 387 118
rect 383 63 387 116
rect 383 61 384 63
rect 386 61 387 63
rect 383 60 387 61
rect 391 110 395 111
rect 391 108 392 110
rect 394 108 395 110
rect 347 37 348 39
rect 350 37 351 39
rect 391 39 395 108
rect 427 63 431 132
rect 567 126 571 127
rect 567 124 568 126
rect 570 124 571 126
rect 471 118 475 119
rect 471 116 472 118
rect 474 116 475 118
rect 427 61 428 63
rect 430 61 431 63
rect 427 60 431 61
rect 435 94 439 95
rect 435 92 436 94
rect 438 92 439 94
rect 391 37 392 39
rect 394 37 395 39
rect 347 36 351 37
rect 379 36 383 37
rect 391 36 395 37
rect 435 39 439 92
rect 471 63 475 116
rect 523 110 527 111
rect 523 108 524 110
rect 526 108 527 110
rect 515 102 519 103
rect 515 100 516 102
rect 518 100 519 102
rect 471 61 472 63
rect 474 61 475 63
rect 471 60 475 61
rect 479 94 483 95
rect 479 92 480 94
rect 482 92 483 94
rect 435 37 436 39
rect 438 37 439 39
rect 435 36 439 37
rect 479 39 483 92
rect 515 63 519 100
rect 515 61 516 63
rect 518 61 519 63
rect 515 60 519 61
rect 479 37 480 39
rect 482 37 483 39
rect 479 36 483 37
rect 523 39 527 108
rect 559 86 563 87
rect 559 84 560 86
rect 562 84 563 86
rect 559 63 563 84
rect 559 61 560 63
rect 562 61 563 63
rect 559 60 563 61
rect 523 37 524 39
rect 526 37 527 39
rect 523 36 527 37
rect 567 39 571 124
rect 611 110 615 111
rect 611 108 612 110
rect 614 108 615 110
rect 603 86 607 87
rect 603 84 604 86
rect 606 84 607 86
rect 603 63 607 84
rect 603 61 604 63
rect 606 61 607 63
rect 603 60 607 61
rect 567 37 568 39
rect 570 37 571 39
rect 567 36 571 37
rect 611 39 615 108
rect 647 102 651 103
rect 647 100 648 102
rect 650 100 651 102
rect 647 63 651 100
rect 647 61 648 63
rect 650 61 651 63
rect 647 60 651 61
rect 655 94 659 95
rect 655 92 656 94
rect 658 92 659 94
rect 611 37 612 39
rect 614 37 615 39
rect 611 36 615 37
rect 655 39 659 92
rect 699 94 703 95
rect 699 92 700 94
rect 702 92 703 94
rect 691 86 695 87
rect 691 84 692 86
rect 694 84 695 86
rect 691 63 695 84
rect 691 61 692 63
rect 694 61 695 63
rect 691 60 695 61
rect 655 37 656 39
rect 658 37 659 39
rect 655 36 659 37
rect 699 39 703 92
rect 730 74 738 77
rect 730 72 733 74
rect 735 72 738 74
rect 730 69 738 72
rect 699 37 700 39
rect 702 37 703 39
rect 699 36 703 37
rect 227 34 228 36
rect 230 34 231 36
rect 227 33 231 34
rect 379 34 380 36
rect 382 34 383 36
rect 183 29 187 30
rect 183 27 184 29
rect 186 27 187 29
rect 183 26 187 27
rect 271 21 275 22
rect 271 19 272 21
rect 274 19 275 21
rect 271 18 275 19
rect 345 21 349 22
rect 345 19 346 21
rect 348 19 349 21
rect 273 -5 277 -4
rect 273 -7 274 -5
rect 276 -7 277 -5
rect 184 -18 188 -17
rect 184 -20 185 -18
rect 187 -20 188 -18
rect 184 -21 188 -20
rect 265 -18 269 -17
rect 265 -20 266 -18
rect 268 -20 269 -18
rect 265 -21 269 -20
rect 152 -27 153 -25
rect 155 -27 156 -25
rect 152 -28 156 -27
rect 201 -26 205 -25
rect 201 -28 202 -26
rect 204 -28 205 -26
rect 201 -29 205 -28
rect 232 -26 236 -25
rect 232 -28 233 -26
rect 235 -28 236 -26
rect 232 -29 236 -28
rect 144 -32 148 -31
rect 144 -34 145 -32
rect 147 -34 148 -32
rect 105 -39 109 -38
rect 105 -41 106 -39
rect 108 -41 109 -39
rect 105 -80 109 -41
rect 105 -82 106 -80
rect 108 -82 109 -80
rect 105 -83 109 -82
rect 128 -103 132 -102
rect 128 -105 129 -103
rect 131 -105 132 -103
rect 128 -106 132 -105
rect 96 -113 97 -111
rect 99 -113 100 -111
rect 96 -114 100 -113
rect 144 -111 148 -34
rect 224 -34 228 -33
rect 224 -36 225 -34
rect 227 -36 228 -34
rect 200 -38 204 -37
rect 200 -40 201 -38
rect 203 -40 204 -38
rect 200 -41 204 -40
rect 209 -94 213 -93
rect 209 -96 210 -94
rect 212 -96 213 -94
rect 209 -97 213 -96
rect 224 -95 228 -36
rect 257 -80 261 -79
rect 257 -82 258 -80
rect 260 -82 261 -80
rect 224 -97 225 -95
rect 227 -97 228 -95
rect 224 -98 228 -97
rect 235 -95 239 -94
rect 235 -97 236 -95
rect 238 -97 239 -95
rect 224 -103 229 -102
rect 224 -105 226 -103
rect 228 -105 229 -103
rect 177 -106 181 -105
rect 177 -108 178 -106
rect 180 -108 181 -106
rect 177 -109 181 -108
rect 208 -106 212 -105
rect 224 -106 229 -105
rect 208 -108 209 -106
rect 211 -108 212 -106
rect 208 -109 212 -108
rect 144 -113 145 -111
rect 147 -113 148 -111
rect 224 -111 228 -110
rect 224 -113 225 -111
rect 227 -113 228 -111
rect 144 -114 148 -113
rect 185 -114 189 -113
rect 185 -116 186 -114
rect 188 -116 189 -114
rect 55 -119 59 -118
rect 55 -121 56 -119
rect 58 -121 59 -119
rect 7 -247 11 -246
rect 7 -249 8 -247
rect 10 -249 11 -247
rect 7 -250 11 -249
rect 55 -255 59 -121
rect 96 -119 100 -118
rect 96 -121 97 -119
rect 99 -121 100 -119
rect 96 -122 100 -121
rect 185 -119 189 -116
rect 185 -121 186 -119
rect 188 -121 189 -119
rect 185 -122 189 -121
rect 66 -134 70 -133
rect 66 -136 67 -134
rect 69 -136 70 -134
rect 66 -242 70 -136
rect 224 -161 228 -113
rect 235 -111 239 -97
rect 257 -98 261 -82
rect 257 -100 258 -98
rect 260 -100 261 -98
rect 257 -102 261 -100
rect 235 -113 236 -111
rect 238 -113 239 -111
rect 235 -114 239 -113
rect 273 -111 277 -7
rect 313 -24 317 -23
rect 313 -26 314 -24
rect 316 -26 317 -24
rect 281 -29 285 -28
rect 281 -31 282 -29
rect 284 -31 285 -29
rect 281 -32 285 -31
rect 313 -75 317 -26
rect 345 -26 349 19
rect 361 21 365 22
rect 361 19 362 21
rect 364 19 365 21
rect 361 18 365 19
rect 370 21 375 22
rect 370 19 371 21
rect 373 19 375 21
rect 345 -28 346 -26
rect 348 -28 349 -26
rect 345 -29 349 -28
rect 362 12 366 14
rect 362 10 363 12
rect 365 10 366 12
rect 321 -38 325 -37
rect 321 -40 322 -38
rect 324 -40 325 -38
rect 321 -41 325 -40
rect 313 -77 314 -75
rect 316 -77 317 -75
rect 313 -78 317 -77
rect 306 -94 310 -93
rect 306 -96 307 -94
rect 309 -96 310 -94
rect 306 -97 310 -96
rect 346 -103 350 -102
rect 346 -105 347 -103
rect 349 -105 350 -103
rect 346 -106 350 -105
rect 273 -113 274 -111
rect 276 -113 277 -111
rect 273 -114 277 -113
rect 362 -111 366 10
rect 370 -25 375 19
rect 379 12 383 34
rect 491 31 495 32
rect 447 30 451 31
rect 447 28 448 30
rect 450 28 451 30
rect 447 27 451 28
rect 483 30 487 31
rect 483 28 484 30
rect 486 28 487 30
rect 491 29 492 31
rect 494 29 495 31
rect 491 28 495 29
rect 523 31 527 32
rect 523 29 524 31
rect 526 29 527 31
rect 404 21 408 22
rect 404 19 405 21
rect 407 19 408 21
rect 404 18 408 19
rect 379 10 380 12
rect 382 10 383 12
rect 379 9 383 10
rect 370 -27 371 -25
rect 373 -27 375 -25
rect 370 -28 375 -27
rect 402 -29 406 -28
rect 402 -31 403 -29
rect 405 -31 406 -29
rect 402 -32 406 -31
rect 427 -94 431 -93
rect 427 -96 428 -94
rect 430 -96 431 -94
rect 427 -97 431 -96
rect 483 -98 487 28
rect 523 -17 527 29
rect 523 -19 524 -17
rect 526 -19 527 -17
rect 523 -20 527 -19
rect 535 30 539 31
rect 535 28 536 30
rect 538 28 539 30
rect 535 -34 539 28
rect 579 21 583 22
rect 579 19 580 21
rect 582 19 583 21
rect 579 18 583 19
rect 612 21 616 22
rect 612 19 613 21
rect 615 19 616 21
rect 612 -17 616 19
rect 612 -19 613 -17
rect 615 -19 616 -17
rect 612 -20 616 -19
rect 628 21 632 22
rect 628 19 629 21
rect 631 19 632 21
rect 628 -25 632 19
rect 742 6 750 10
rect 742 4 745 6
rect 747 4 750 6
rect 742 0 750 4
rect 628 -27 629 -25
rect 631 -27 632 -25
rect 628 -28 632 -27
rect 535 -36 536 -34
rect 538 -36 539 -34
rect 535 -37 539 -36
rect 571 -33 575 -32
rect 571 -35 572 -33
rect 574 -35 575 -33
rect 491 -39 495 -37
rect 491 -41 492 -39
rect 494 -41 495 -39
rect 491 -51 495 -41
rect 491 -53 492 -51
rect 494 -53 495 -51
rect 491 -54 495 -53
rect 552 -51 556 -50
rect 552 -53 553 -51
rect 555 -53 556 -51
rect 483 -100 484 -98
rect 486 -100 487 -98
rect 483 -101 487 -100
rect 491 -83 495 -82
rect 491 -85 492 -83
rect 494 -85 495 -83
rect 443 -103 447 -102
rect 443 -105 444 -103
rect 446 -105 447 -103
rect 395 -106 399 -105
rect 395 -108 396 -106
rect 398 -108 399 -106
rect 395 -109 399 -108
rect 426 -106 430 -105
rect 443 -106 447 -105
rect 426 -108 427 -106
rect 429 -108 430 -106
rect 426 -109 430 -108
rect 491 -111 495 -85
rect 524 -94 528 -93
rect 524 -96 525 -94
rect 527 -96 528 -94
rect 524 -97 528 -96
rect 362 -113 363 -111
rect 365 -113 366 -111
rect 362 -114 366 -113
rect 403 -112 407 -111
rect 403 -114 404 -112
rect 406 -114 407 -112
rect 491 -113 492 -111
rect 494 -113 495 -111
rect 491 -114 495 -113
rect 552 -111 556 -53
rect 571 -83 575 -35
rect 571 -85 572 -83
rect 574 -85 575 -83
rect 571 -86 575 -85
rect 580 -39 584 -37
rect 580 -41 581 -39
rect 583 -41 584 -39
rect 564 -103 568 -102
rect 564 -105 565 -103
rect 567 -105 568 -103
rect 564 -106 568 -105
rect 552 -113 553 -111
rect 555 -113 556 -111
rect 552 -114 556 -113
rect 560 -111 564 -110
rect 560 -113 561 -111
rect 563 -113 564 -111
rect 314 -117 318 -116
rect 279 -119 283 -118
rect 279 -121 280 -119
rect 282 -121 283 -119
rect 279 -150 283 -121
rect 314 -119 315 -117
rect 317 -119 318 -117
rect 314 -149 318 -119
rect 403 -134 407 -114
rect 403 -136 404 -134
rect 406 -136 407 -134
rect 403 -137 407 -136
rect 279 -152 280 -150
rect 282 -152 283 -150
rect 279 -153 283 -152
rect 292 -150 296 -149
rect 292 -152 293 -150
rect 295 -152 296 -150
rect 314 -151 315 -149
rect 317 -151 318 -149
rect 314 -152 318 -151
rect 416 -149 420 -148
rect 416 -151 417 -149
rect 419 -151 420 -149
rect 224 -163 225 -161
rect 227 -163 228 -161
rect 224 -164 228 -163
rect 241 -170 245 -169
rect 241 -172 242 -170
rect 244 -172 245 -170
rect 241 -173 245 -172
rect 283 -170 287 -169
rect 283 -172 284 -170
rect 286 -172 287 -170
rect 283 -173 287 -172
rect 264 -177 268 -176
rect 264 -179 265 -177
rect 267 -179 268 -177
rect 240 -182 244 -181
rect 240 -184 241 -182
rect 243 -184 244 -182
rect 240 -185 244 -184
rect 155 -208 159 -207
rect 155 -210 156 -208
rect 158 -210 159 -208
rect 88 -238 92 -237
rect 88 -240 89 -238
rect 91 -240 92 -238
rect 88 -241 92 -240
rect 66 -244 67 -242
rect 69 -244 70 -242
rect 66 -245 70 -244
rect 139 -247 143 -246
rect 139 -249 140 -247
rect 142 -249 143 -247
rect 139 -250 143 -249
rect 55 -257 56 -255
rect 58 -257 59 -255
rect 55 -258 59 -257
rect 155 -255 159 -210
rect 264 -208 268 -179
rect 264 -210 265 -208
rect 267 -210 268 -208
rect 264 -211 268 -210
rect 279 -190 283 -187
rect 279 -192 280 -190
rect 282 -192 283 -190
rect 231 -238 235 -237
rect 231 -240 232 -238
rect 234 -240 235 -238
rect 231 -241 235 -240
rect 279 -242 283 -192
rect 292 -190 296 -152
rect 316 -161 320 -160
rect 316 -163 317 -161
rect 319 -163 320 -161
rect 316 -164 320 -163
rect 416 -161 420 -151
rect 416 -163 417 -161
rect 419 -163 420 -161
rect 416 -164 420 -163
rect 560 -162 564 -113
rect 580 -111 584 -41
rect 727 -66 739 -62
rect 727 -68 732 -66
rect 734 -68 739 -66
rect 727 -71 739 -68
rect 660 -75 664 -74
rect 660 -77 661 -75
rect 663 -77 664 -75
rect 645 -94 649 -93
rect 645 -96 646 -94
rect 648 -96 649 -94
rect 645 -97 649 -96
rect 613 -106 617 -105
rect 613 -108 614 -106
rect 616 -108 617 -106
rect 613 -109 617 -108
rect 644 -106 648 -105
rect 644 -108 645 -106
rect 647 -108 648 -106
rect 644 -109 648 -108
rect 580 -113 581 -111
rect 583 -113 584 -111
rect 580 -114 584 -113
rect 621 -115 625 -114
rect 621 -117 622 -115
rect 624 -117 625 -115
rect 621 -118 625 -117
rect 560 -164 561 -162
rect 563 -164 564 -162
rect 660 -161 664 -77
rect 660 -163 661 -161
rect 663 -163 664 -161
rect 660 -164 664 -163
rect 668 -115 672 -114
rect 668 -117 669 -115
rect 671 -117 672 -115
rect 560 -165 564 -164
rect 485 -170 489 -169
rect 485 -172 486 -170
rect 488 -172 489 -170
rect 332 -173 336 -172
rect 332 -175 333 -173
rect 335 -175 336 -173
rect 332 -176 336 -175
rect 464 -173 468 -172
rect 485 -173 489 -172
rect 527 -170 531 -169
rect 527 -172 528 -170
rect 530 -172 531 -170
rect 527 -173 531 -172
rect 576 -173 580 -172
rect 464 -175 465 -173
rect 467 -175 468 -173
rect 464 -176 468 -175
rect 576 -175 577 -173
rect 579 -175 580 -173
rect 576 -176 580 -175
rect 433 -178 437 -177
rect 433 -180 434 -178
rect 436 -180 437 -178
rect 383 -182 387 -181
rect 383 -184 384 -182
rect 386 -184 387 -182
rect 383 -185 387 -184
rect 292 -192 293 -190
rect 295 -192 296 -190
rect 292 -193 296 -192
rect 433 -194 437 -180
rect 668 -178 672 -117
rect 747 -138 755 -134
rect 747 -140 750 -138
rect 752 -140 755 -138
rect 747 -144 755 -140
rect 708 -173 712 -172
rect 708 -175 709 -173
rect 711 -175 712 -173
rect 708 -176 712 -175
rect 668 -180 669 -178
rect 671 -180 672 -178
rect 668 -181 672 -180
rect 484 -182 488 -181
rect 484 -184 485 -182
rect 487 -184 488 -182
rect 484 -185 488 -184
rect 627 -182 631 -181
rect 627 -184 628 -182
rect 630 -184 631 -182
rect 627 -185 631 -184
rect 433 -196 434 -194
rect 436 -196 437 -194
rect 433 -197 437 -196
rect 499 -194 503 -193
rect 499 -196 500 -194
rect 502 -196 503 -194
rect 499 -197 503 -196
rect 734 -206 742 -203
rect 734 -208 737 -206
rect 739 -208 742 -206
rect 734 -211 742 -208
rect 329 -238 333 -237
rect 329 -240 330 -238
rect 332 -240 333 -238
rect 329 -241 333 -240
rect 472 -238 476 -237
rect 472 -240 473 -238
rect 475 -240 476 -238
rect 472 -241 476 -240
rect 279 -244 280 -242
rect 282 -244 283 -242
rect 279 -245 283 -244
rect 248 -247 252 -246
rect 248 -249 249 -247
rect 251 -249 252 -247
rect 188 -250 192 -249
rect 188 -252 189 -250
rect 191 -252 192 -250
rect 188 -253 192 -252
rect 230 -250 234 -249
rect 248 -250 252 -249
rect 380 -247 384 -246
rect 380 -249 381 -247
rect 383 -249 384 -247
rect 380 -250 384 -249
rect 429 -250 433 -249
rect 230 -252 231 -250
rect 233 -252 234 -250
rect 230 -253 234 -252
rect 429 -252 430 -250
rect 432 -252 433 -250
rect 429 -253 433 -252
rect 471 -250 475 -249
rect 471 -252 472 -250
rect 474 -252 475 -250
rect 471 -253 475 -252
rect 155 -257 156 -255
rect 158 -257 159 -255
rect 155 -258 159 -257
rect 207 -258 211 -257
rect 207 -260 208 -258
rect 210 -260 211 -258
rect 207 -261 211 -260
rect 296 -258 300 -257
rect 296 -260 297 -258
rect 299 -260 300 -258
rect 296 -261 300 -260
rect 396 -259 400 -258
rect 396 -261 397 -259
rect 399 -261 400 -259
rect -1 -282 0 -280
rect 2 -282 3 -280
rect -1 -283 3 -282
rect 396 -280 400 -261
rect 396 -282 397 -280
rect 399 -282 400 -280
rect 396 -283 400 -282
rect 715 -278 726 -275
rect 715 -280 719 -278
rect 721 -280 726 -278
rect 715 -283 726 -280
<< alu3 >>
rect -22 74 -15 77
rect -22 72 -19 74
rect -17 72 -15 74
rect -22 69 -15 72
rect 730 74 738 77
rect 730 72 733 74
rect 735 72 738 74
rect 730 69 738 72
rect 152 55 319 56
rect 152 53 153 55
rect 155 53 316 55
rect 318 53 319 55
rect 152 52 319 53
rect 47 38 143 39
rect 47 36 48 38
rect 50 36 140 38
rect 142 36 143 38
rect 47 35 143 36
rect 227 36 383 37
rect 227 34 228 36
rect 230 34 380 36
rect 382 34 383 36
rect 227 33 383 34
rect -1 31 11 32
rect 491 31 527 32
rect -1 29 0 31
rect 2 29 8 31
rect 10 29 11 31
rect 447 30 487 31
rect -1 28 11 29
rect 63 29 187 30
rect 63 27 64 29
rect 66 27 184 29
rect 186 27 187 29
rect 447 28 448 30
rect 450 28 484 30
rect 486 28 487 30
rect 491 29 492 31
rect 494 29 524 31
rect 526 29 527 31
rect 491 28 527 29
rect 447 27 487 28
rect 63 26 187 27
rect 136 21 275 22
rect 136 19 137 21
rect 139 19 272 21
rect 274 19 275 21
rect 136 18 275 19
rect 345 21 365 22
rect 345 19 346 21
rect 348 19 362 21
rect 364 19 365 21
rect 345 18 365 19
rect 370 21 409 22
rect 370 19 371 21
rect 373 19 405 21
rect 407 19 409 21
rect 370 18 409 19
rect 579 21 616 22
rect 579 19 580 21
rect 582 19 613 21
rect 615 19 616 21
rect 579 18 616 19
rect -24 6 -12 13
rect 362 12 383 13
rect 362 10 363 12
rect 365 10 380 12
rect 382 10 383 12
rect 362 9 383 10
rect -24 4 -19 6
rect -17 4 -12 6
rect -24 -3 -12 4
rect 742 6 750 10
rect 742 4 745 6
rect 747 4 750 6
rect 742 0 750 4
rect 88 -5 277 -4
rect 88 -7 89 -5
rect 91 -7 274 -5
rect 276 -7 277 -5
rect 88 -8 277 -7
rect 184 -18 269 -17
rect 184 -20 185 -18
rect 187 -20 266 -18
rect 268 -20 269 -18
rect 184 -21 269 -20
rect 201 -26 236 -25
rect 201 -28 202 -26
rect 204 -28 233 -26
rect 235 -28 236 -26
rect 201 -29 236 -28
rect 281 -29 406 -28
rect 281 -31 282 -29
rect 284 -31 403 -29
rect 405 -31 406 -29
rect 14 -32 148 -31
rect 281 -32 406 -31
rect 14 -34 15 -32
rect 17 -34 145 -32
rect 147 -34 148 -32
rect 14 -35 148 -34
rect 200 -38 325 -37
rect 200 -40 201 -38
rect 203 -40 322 -38
rect 324 -40 325 -38
rect 200 -41 325 -40
rect 491 -51 556 -50
rect 491 -53 492 -51
rect 494 -53 553 -51
rect 555 -53 556 -51
rect 491 -54 556 -53
rect -21 -66 -15 -63
rect -21 -68 -19 -66
rect -17 -68 -15 -66
rect -21 -71 -15 -68
rect 727 -66 739 -62
rect 727 -68 732 -66
rect 734 -68 739 -66
rect 727 -71 739 -68
rect 313 -75 664 -74
rect 313 -77 314 -75
rect 316 -77 661 -75
rect 663 -77 664 -75
rect 313 -78 664 -77
rect 105 -80 261 -79
rect 105 -82 106 -80
rect 108 -82 258 -80
rect 260 -82 261 -80
rect 105 -83 261 -82
rect 491 -83 575 -82
rect 491 -85 492 -83
rect 494 -85 572 -83
rect 574 -85 575 -83
rect 491 -86 575 -85
rect 88 -94 213 -93
rect 306 -94 431 -93
rect 88 -96 89 -94
rect 91 -96 210 -94
rect 212 -96 213 -94
rect 88 -97 213 -96
rect 224 -95 239 -94
rect 224 -97 225 -95
rect 227 -97 236 -95
rect 238 -97 239 -95
rect 306 -96 307 -94
rect 309 -96 428 -94
rect 430 -96 431 -94
rect 306 -97 431 -96
rect 524 -94 649 -93
rect 524 -96 525 -94
rect 527 -96 646 -94
rect 648 -96 649 -94
rect 524 -97 649 -96
rect 224 -98 239 -97
rect 7 -103 132 -102
rect 7 -105 8 -103
rect 10 -105 129 -103
rect 131 -105 132 -103
rect 225 -103 350 -102
rect 225 -105 226 -103
rect 228 -105 347 -103
rect 349 -105 350 -103
rect 443 -103 568 -102
rect 443 -105 444 -103
rect 446 -105 565 -103
rect 567 -105 568 -103
rect 7 -106 132 -105
rect 177 -106 212 -105
rect 225 -106 350 -105
rect 395 -106 430 -105
rect 443 -106 568 -105
rect 613 -106 648 -105
rect 177 -108 178 -106
rect 180 -108 209 -106
rect 211 -108 212 -106
rect 177 -109 212 -108
rect 395 -108 396 -106
rect 398 -108 427 -106
rect 429 -108 430 -106
rect 395 -109 430 -108
rect 613 -108 614 -106
rect 616 -108 645 -106
rect 647 -108 648 -106
rect 613 -109 648 -108
rect 55 -111 100 -110
rect 55 -113 56 -111
rect 58 -113 97 -111
rect 99 -113 100 -111
rect 55 -114 100 -113
rect 224 -111 239 -110
rect 224 -113 225 -111
rect 227 -113 236 -111
rect 238 -113 239 -111
rect 224 -114 239 -113
rect 552 -111 564 -110
rect 552 -113 553 -111
rect 555 -113 561 -111
rect 563 -113 564 -111
rect 552 -114 564 -113
rect 621 -115 672 -114
rect 621 -117 622 -115
rect 624 -117 669 -115
rect 671 -117 672 -115
rect 621 -118 672 -117
rect 55 -119 100 -118
rect 55 -121 56 -119
rect 58 -121 97 -119
rect 99 -121 100 -119
rect 55 -122 100 -121
rect 185 -119 283 -118
rect 185 -121 186 -119
rect 188 -121 280 -119
rect 282 -121 283 -119
rect 185 -122 283 -121
rect -30 -134 -24 -131
rect -30 -136 -28 -134
rect -26 -136 -24 -134
rect -30 -139 -24 -136
rect 66 -134 407 -133
rect 66 -136 67 -134
rect 69 -136 404 -134
rect 406 -136 407 -134
rect 66 -137 407 -136
rect 747 -138 755 -134
rect 747 -140 750 -138
rect 752 -140 755 -138
rect 747 -144 755 -140
rect 314 -149 420 -148
rect 279 -150 296 -149
rect 279 -152 280 -150
rect 282 -152 293 -150
rect 295 -152 296 -150
rect 314 -151 315 -149
rect 317 -151 417 -149
rect 419 -151 420 -149
rect 314 -152 420 -151
rect 279 -153 296 -152
rect 224 -161 320 -160
rect 224 -163 225 -161
rect 227 -163 317 -161
rect 319 -163 320 -161
rect 224 -164 320 -163
rect 241 -170 287 -169
rect 241 -172 242 -170
rect 244 -172 284 -170
rect 286 -172 287 -170
rect 485 -170 531 -169
rect 485 -172 486 -170
rect 488 -172 528 -170
rect 530 -172 531 -170
rect 241 -173 287 -172
rect 332 -173 468 -172
rect 485 -173 531 -172
rect 576 -173 712 -172
rect 332 -175 333 -173
rect 335 -175 465 -173
rect 467 -175 468 -173
rect 332 -176 468 -175
rect 576 -175 577 -173
rect 579 -175 709 -173
rect 711 -175 712 -173
rect 576 -176 712 -175
rect 240 -182 387 -181
rect 240 -184 241 -182
rect 243 -184 384 -182
rect 386 -184 387 -182
rect 240 -185 387 -184
rect 484 -182 631 -181
rect 484 -184 485 -182
rect 487 -184 628 -182
rect 630 -184 631 -182
rect 484 -185 631 -184
rect 279 -190 296 -189
rect 279 -192 280 -190
rect 282 -192 293 -190
rect 295 -192 296 -190
rect 279 -193 296 -192
rect 433 -194 503 -193
rect 433 -196 434 -194
rect 436 -196 500 -194
rect 502 -196 503 -194
rect 433 -197 503 -196
rect 734 -206 742 -203
rect -22 -210 -15 -207
rect -22 -212 -20 -210
rect -18 -212 -15 -210
rect 155 -208 268 -207
rect 155 -210 156 -208
rect 158 -210 265 -208
rect 267 -210 268 -208
rect 155 -211 268 -210
rect 734 -208 737 -206
rect 739 -208 742 -206
rect 734 -211 742 -208
rect -22 -215 -15 -212
rect 88 -238 235 -237
rect 88 -240 89 -238
rect 91 -240 232 -238
rect 234 -240 235 -238
rect 88 -241 235 -240
rect 329 -238 476 -237
rect 329 -240 330 -238
rect 332 -240 473 -238
rect 475 -240 476 -238
rect 329 -241 476 -240
rect 7 -247 143 -246
rect 7 -249 8 -247
rect 10 -249 140 -247
rect 142 -249 143 -247
rect 248 -247 384 -246
rect 248 -249 249 -247
rect 251 -249 381 -247
rect 383 -249 384 -247
rect 7 -250 143 -249
rect 188 -250 234 -249
rect 248 -250 384 -249
rect 429 -250 475 -249
rect 188 -252 189 -250
rect 191 -252 231 -250
rect 233 -252 234 -250
rect 188 -253 234 -252
rect 429 -252 430 -250
rect 432 -252 472 -250
rect 474 -252 475 -250
rect 429 -253 475 -252
rect 207 -258 300 -257
rect 207 -260 208 -258
rect 210 -260 297 -258
rect 299 -260 300 -258
rect 207 -261 300 -260
rect -33 -278 -27 -275
rect -33 -280 -31 -278
rect -29 -280 -27 -278
rect 715 -278 726 -275
rect -33 -282 -27 -280
rect -1 -280 400 -279
rect -1 -282 0 -280
rect 2 -282 397 -280
rect 399 -282 400 -280
rect -1 -283 400 -282
rect 715 -280 719 -278
rect 721 -280 726 -278
rect 715 -283 726 -280
<< alu4 >>
rect -22 74 -15 77
rect -22 72 -19 74
rect -17 72 -15 74
rect -22 69 -15 72
rect 730 74 738 77
rect 730 72 733 74
rect 735 72 738 74
rect 730 69 738 72
rect -24 6 -12 13
rect -24 4 -19 6
rect -17 4 -12 6
rect -24 -3 -12 4
rect 742 6 750 10
rect 742 4 745 6
rect 747 4 750 6
rect 742 0 750 4
rect -21 -66 -15 -63
rect -21 -68 -19 -66
rect -17 -68 -15 -66
rect -21 -71 -15 -68
rect 727 -66 739 -62
rect 727 -68 732 -66
rect 734 -68 739 -66
rect 727 -71 739 -68
rect -30 -134 -24 -131
rect -30 -136 -28 -134
rect -26 -136 -24 -134
rect -30 -139 -24 -136
rect 747 -138 755 -134
rect 747 -140 750 -138
rect 752 -140 755 -138
rect 747 -144 755 -140
rect 734 -206 742 -203
rect -22 -210 -15 -207
rect -22 -212 -20 -210
rect -18 -212 -15 -210
rect 734 -208 737 -206
rect 739 -208 742 -206
rect 734 -211 742 -208
rect -22 -215 -15 -212
rect -33 -278 -27 -275
rect -33 -280 -31 -278
rect -29 -280 -27 -278
rect -33 -282 -27 -280
rect 715 -278 726 -275
rect 715 -280 719 -278
rect 721 -280 726 -278
rect 715 -283 726 -280
<< alu5 >>
rect -111 222 834 226
rect -111 218 -107 222
rect -103 218 826 222
rect 830 218 834 222
rect -111 214 834 218
rect -59 191 780 195
rect -59 187 -55 191
rect -51 187 772 191
rect 776 187 780 191
rect -59 183 780 187
rect -111 75 -15 77
rect -111 71 -107 75
rect -103 74 -15 75
rect -103 72 -19 74
rect -17 72 -15 74
rect -103 71 -15 72
rect -111 69 -15 71
rect 730 75 834 77
rect 730 74 826 75
rect 730 72 733 74
rect 735 72 826 74
rect 730 71 826 72
rect 830 71 834 75
rect 730 69 834 71
rect -59 8 -12 13
rect 768 10 780 12
rect -59 4 -55 8
rect -51 6 -12 8
rect -51 4 -19 6
rect -17 4 -12 6
rect -59 -3 -12 4
rect 742 8 780 10
rect 742 6 772 8
rect 742 4 745 6
rect 747 4 772 6
rect 776 4 780 8
rect 742 0 780 4
rect -111 -65 -15 -63
rect -111 -69 -107 -65
rect -103 -66 -15 -65
rect -103 -68 -19 -66
rect -17 -68 -15 -66
rect -103 -69 -15 -68
rect -111 -71 -15 -69
rect 727 -65 834 -62
rect 727 -66 826 -65
rect 727 -68 732 -66
rect 734 -68 826 -66
rect 727 -69 826 -68
rect 830 -69 834 -65
rect 727 -71 834 -69
rect -59 -133 -24 -131
rect -59 -137 -55 -133
rect -51 -134 -24 -133
rect 768 -134 780 -132
rect -51 -136 -28 -134
rect -26 -136 -24 -134
rect -51 -137 -24 -136
rect -59 -139 -24 -137
rect 747 -136 780 -134
rect 747 -138 772 -136
rect 747 -140 750 -138
rect 752 -140 772 -138
rect 776 -140 780 -136
rect 747 -144 780 -140
rect -111 -207 -99 -203
rect 734 -205 834 -203
rect 734 -206 826 -205
rect -111 -209 -15 -207
rect -111 -213 -107 -209
rect -103 -210 -15 -209
rect -103 -212 -20 -210
rect -18 -212 -15 -210
rect 734 -208 737 -206
rect 739 -208 826 -206
rect 734 -209 826 -208
rect 830 -209 834 -205
rect 734 -211 834 -209
rect -103 -213 -15 -212
rect -111 -215 -15 -213
rect -59 -275 -45 -274
rect 768 -275 780 -272
rect -59 -276 -27 -275
rect -59 -280 -55 -276
rect -51 -278 -27 -276
rect -51 -280 -31 -278
rect -29 -280 -27 -278
rect -59 -282 -27 -280
rect 715 -277 780 -275
rect 715 -278 772 -277
rect 715 -280 719 -278
rect 721 -280 772 -278
rect 715 -281 772 -280
rect 776 -281 780 -277
rect 715 -283 780 -281
rect 768 -284 780 -283
rect -59 -329 780 -325
rect -59 -333 -55 -329
rect -51 -333 772 -329
rect 776 -333 780 -329
rect -59 -337 780 -333
rect -111 -357 834 -353
rect -111 -361 -107 -357
rect -103 -361 826 -357
rect 830 -361 834 -357
rect -111 -365 834 -361
<< alu6 >>
rect -111 222 -99 226
rect -111 218 -107 222
rect -103 218 -99 222
rect -111 75 -99 218
rect 822 222 834 226
rect 822 218 826 222
rect 830 218 834 222
rect -111 71 -107 75
rect -103 71 -99 75
rect -111 -65 -99 71
rect -111 -69 -107 -65
rect -103 -69 -99 -65
rect -111 -209 -99 -69
rect -111 -213 -107 -209
rect -103 -213 -99 -209
rect -111 -357 -99 -213
rect -59 191 -47 195
rect -59 187 -55 191
rect -51 187 -47 191
rect -59 8 -47 187
rect -59 4 -55 8
rect -51 4 -47 8
rect -59 -133 -47 4
rect -59 -137 -55 -133
rect -51 -137 -47 -133
rect -59 -276 -47 -137
rect -59 -280 -55 -276
rect -51 -280 -47 -276
rect -59 -329 -47 -280
rect -59 -333 -55 -329
rect -51 -333 -47 -329
rect -59 -337 -47 -333
rect 768 191 780 195
rect 768 187 772 191
rect 776 187 780 191
rect 768 8 780 187
rect 768 4 772 8
rect 776 4 780 8
rect 768 -136 780 4
rect 768 -140 772 -136
rect 776 -140 780 -136
rect 768 -277 780 -140
rect 768 -281 772 -277
rect 776 -281 780 -277
rect 768 -329 780 -281
rect 768 -333 772 -329
rect 776 -333 780 -329
rect 768 -337 780 -333
rect 822 75 834 218
rect 822 71 826 75
rect 830 71 834 75
rect 822 -65 834 71
rect 822 -69 826 -65
rect 830 -69 834 -65
rect 822 -205 834 -69
rect 822 -209 826 -205
rect 830 -209 834 -205
rect -111 -361 -107 -357
rect -103 -361 -99 -357
rect -111 -365 -99 -361
rect 822 -357 834 -209
rect 822 -361 826 -357
rect 830 -361 834 -357
rect 822 -365 834 -361
<< ptie >>
rect 8 12 14 14
rect 8 10 10 12
rect 12 10 14 12
rect 8 8 14 10
rect 52 12 58 14
rect 52 10 54 12
rect 56 10 58 12
rect 52 8 58 10
rect 96 12 102 14
rect 96 10 98 12
rect 100 10 102 12
rect 96 8 102 10
rect 140 12 146 14
rect 140 10 142 12
rect 144 10 146 12
rect 140 8 146 10
rect 184 12 190 14
rect 184 10 186 12
rect 188 10 190 12
rect 184 8 190 10
rect 228 12 234 14
rect 228 10 230 12
rect 232 10 234 12
rect 228 8 234 10
rect 272 12 278 14
rect 272 10 274 12
rect 276 10 278 12
rect 272 8 278 10
rect 316 12 322 14
rect 316 10 318 12
rect 320 10 322 12
rect 316 8 322 10
rect 360 12 366 14
rect 360 10 362 12
rect 364 10 366 12
rect 360 8 366 10
rect 404 12 410 14
rect 404 10 406 12
rect 408 10 410 12
rect 404 8 410 10
rect 448 12 454 14
rect 448 10 450 12
rect 452 10 454 12
rect 448 8 454 10
rect 492 12 498 14
rect 492 10 494 12
rect 496 10 498 12
rect 492 8 498 10
rect 536 12 542 14
rect 536 10 538 12
rect 540 10 542 12
rect 536 8 542 10
rect 580 12 586 14
rect 580 10 582 12
rect 584 10 586 12
rect 580 8 586 10
rect 624 12 630 14
rect 624 10 626 12
rect 628 10 630 12
rect 624 8 630 10
rect 668 12 674 14
rect 668 10 670 12
rect 672 10 674 12
rect 668 8 674 10
rect 193 0 227 2
rect 193 -2 195 0
rect 197 -2 223 0
rect 225 -2 227 0
rect 193 -4 227 -2
rect 186 -132 220 -130
rect 186 -134 188 -132
rect 190 -134 216 -132
rect 218 -134 220 -132
rect 186 -136 220 -134
rect 404 -132 438 -130
rect 404 -134 406 -132
rect 408 -134 434 -132
rect 436 -134 438 -132
rect 404 -136 438 -134
rect 622 -132 656 -130
rect 622 -134 624 -132
rect 626 -134 652 -132
rect 654 -134 656 -132
rect 622 -136 656 -134
rect 233 -144 267 -142
rect 233 -146 235 -144
rect 237 -146 263 -144
rect 265 -146 267 -144
rect 233 -148 267 -146
rect 477 -144 511 -142
rect 477 -146 479 -144
rect 481 -146 507 -144
rect 509 -146 511 -144
rect 477 -148 511 -146
rect 208 -276 242 -274
rect 208 -278 210 -276
rect 212 -278 238 -276
rect 240 -278 242 -276
rect 208 -280 242 -278
rect 449 -276 483 -274
rect 449 -278 451 -276
rect 453 -278 479 -276
rect 481 -278 483 -276
rect 449 -280 483 -278
<< ntie >>
rect 8 72 42 74
rect 8 70 10 72
rect 12 70 24 72
rect 26 70 38 72
rect 40 70 42 72
rect 8 68 42 70
rect 52 72 86 74
rect 52 70 54 72
rect 56 70 68 72
rect 70 70 82 72
rect 84 70 86 72
rect 52 68 86 70
rect 96 72 130 74
rect 96 70 98 72
rect 100 70 112 72
rect 114 70 126 72
rect 128 70 130 72
rect 96 68 130 70
rect 140 72 174 74
rect 140 70 142 72
rect 144 70 156 72
rect 158 70 170 72
rect 172 70 174 72
rect 140 68 174 70
rect 184 72 218 74
rect 184 70 186 72
rect 188 70 200 72
rect 202 70 214 72
rect 216 70 218 72
rect 184 68 218 70
rect 228 72 262 74
rect 228 70 230 72
rect 232 70 244 72
rect 246 70 258 72
rect 260 70 262 72
rect 228 68 262 70
rect 272 72 306 74
rect 272 70 274 72
rect 276 70 288 72
rect 290 70 302 72
rect 304 70 306 72
rect 272 68 306 70
rect 316 72 350 74
rect 316 70 318 72
rect 320 70 332 72
rect 334 70 346 72
rect 348 70 350 72
rect 316 68 350 70
rect 360 72 394 74
rect 360 70 362 72
rect 364 70 376 72
rect 378 70 390 72
rect 392 70 394 72
rect 360 68 394 70
rect 404 72 438 74
rect 404 70 406 72
rect 408 70 420 72
rect 422 70 434 72
rect 436 70 438 72
rect 404 68 438 70
rect 448 72 482 74
rect 448 70 450 72
rect 452 70 464 72
rect 466 70 478 72
rect 480 70 482 72
rect 448 68 482 70
rect 492 72 526 74
rect 492 70 494 72
rect 496 70 508 72
rect 510 70 522 72
rect 524 70 526 72
rect 492 68 526 70
rect 536 72 570 74
rect 536 70 538 72
rect 540 70 552 72
rect 554 70 566 72
rect 568 70 570 72
rect 536 68 570 70
rect 580 72 614 74
rect 580 70 582 72
rect 584 70 596 72
rect 598 70 610 72
rect 612 70 614 72
rect 580 68 614 70
rect 624 72 658 74
rect 624 70 626 72
rect 628 70 640 72
rect 642 70 654 72
rect 656 70 658 72
rect 624 68 658 70
rect 668 72 702 74
rect 668 70 670 72
rect 672 70 684 72
rect 686 70 698 72
rect 700 70 702 72
rect 668 68 702 70
rect 221 -60 227 -58
rect 221 -62 223 -60
rect 225 -62 227 -60
rect 221 -64 227 -62
rect 186 -72 192 -70
rect 186 -74 188 -72
rect 190 -74 192 -72
rect 186 -76 192 -74
rect 404 -72 410 -70
rect 404 -74 406 -72
rect 408 -74 410 -72
rect 404 -76 410 -74
rect 622 -72 628 -70
rect 622 -74 624 -72
rect 626 -74 628 -72
rect 622 -76 628 -74
rect 261 -204 267 -202
rect 261 -206 263 -204
rect 265 -206 267 -204
rect 261 -208 267 -206
rect 505 -204 511 -202
rect 505 -206 507 -204
rect 509 -206 511 -204
rect 505 -208 511 -206
rect 208 -216 214 -214
rect 208 -218 210 -216
rect 212 -218 214 -216
rect 208 -220 214 -218
rect 449 -216 455 -214
rect 449 -218 451 -216
rect 453 -218 455 -216
rect 449 -220 455 -218
<< nmos >>
rect 14 20 16 26
rect 26 14 28 23
rect 33 14 35 23
rect 58 20 60 26
rect 70 14 72 23
rect 77 14 79 23
rect 102 20 104 26
rect 114 14 116 23
rect 121 14 123 23
rect 146 20 148 26
rect 158 14 160 23
rect 165 14 167 23
rect 190 20 192 26
rect 202 14 204 23
rect 209 14 211 23
rect 234 20 236 26
rect 246 14 248 23
rect 253 14 255 23
rect 278 20 280 26
rect 290 14 292 23
rect 297 14 299 23
rect 322 20 324 26
rect 334 14 336 23
rect 341 14 343 23
rect 366 20 368 26
rect 378 14 380 23
rect 385 14 387 23
rect 410 20 412 26
rect 422 14 424 23
rect 429 14 431 23
rect 454 20 456 26
rect 466 14 468 23
rect 473 14 475 23
rect 498 20 500 26
rect 510 14 512 23
rect 517 14 519 23
rect 542 20 544 26
rect 554 14 556 23
rect 561 14 563 23
rect 586 20 588 26
rect 598 14 600 23
rect 605 14 607 23
rect 630 20 632 26
rect 642 14 644 23
rect 649 14 651 23
rect 674 20 676 26
rect 686 14 688 23
rect 693 14 695 23
rect 22 -15 24 -1
rect 33 -21 35 -1
rect 40 -21 42 -1
rect 60 -21 62 -7
rect 70 -21 72 -7
rect 80 -14 82 -4
rect 90 -14 92 -1
rect 111 -15 113 -1
rect 122 -21 124 -1
rect 129 -21 131 -1
rect 149 -21 151 -7
rect 159 -21 161 -7
rect 169 -14 171 -4
rect 179 -14 181 -1
rect 199 -16 201 -10
rect 209 -16 211 -10
rect 219 -16 221 -10
rect 240 -15 242 -1
rect 251 -21 253 -1
rect 258 -21 260 -1
rect 278 -21 280 -7
rect 288 -21 290 -7
rect 298 -14 300 -4
rect 308 -14 310 -1
rect 329 -15 331 -1
rect 340 -21 342 -1
rect 347 -21 349 -1
rect 367 -21 369 -7
rect 377 -21 379 -7
rect 387 -14 389 -4
rect 397 -14 399 -1
rect 498 -15 500 -1
rect 509 -21 511 -1
rect 516 -21 518 -1
rect 536 -21 538 -7
rect 546 -21 548 -7
rect 556 -14 558 -4
rect 566 -14 568 -1
rect 587 -15 589 -1
rect 598 -21 600 -1
rect 605 -21 607 -1
rect 625 -21 627 -7
rect 635 -21 637 -7
rect 645 -14 647 -4
rect 655 -14 657 -1
rect 14 -133 16 -120
rect 24 -130 26 -120
rect 34 -127 36 -113
rect 44 -127 46 -113
rect 64 -133 66 -113
rect 71 -133 73 -113
rect 82 -133 84 -119
rect 103 -133 105 -120
rect 113 -130 115 -120
rect 123 -127 125 -113
rect 133 -127 135 -113
rect 153 -133 155 -113
rect 160 -133 162 -113
rect 171 -133 173 -119
rect 192 -124 194 -118
rect 202 -124 204 -118
rect 212 -124 214 -118
rect 232 -133 234 -120
rect 242 -130 244 -120
rect 252 -127 254 -113
rect 262 -127 264 -113
rect 282 -133 284 -113
rect 289 -133 291 -113
rect 300 -133 302 -119
rect 321 -133 323 -120
rect 331 -130 333 -120
rect 341 -127 343 -113
rect 351 -127 353 -113
rect 371 -133 373 -113
rect 378 -133 380 -113
rect 389 -133 391 -119
rect 410 -124 412 -118
rect 420 -124 422 -118
rect 430 -124 432 -118
rect 450 -133 452 -120
rect 460 -130 462 -120
rect 470 -127 472 -113
rect 480 -127 482 -113
rect 500 -133 502 -113
rect 507 -133 509 -113
rect 518 -133 520 -119
rect 539 -133 541 -120
rect 549 -130 551 -120
rect 559 -127 561 -113
rect 569 -127 571 -113
rect 589 -133 591 -113
rect 596 -133 598 -113
rect 607 -133 609 -119
rect 628 -124 630 -118
rect 638 -124 640 -118
rect 648 -124 650 -118
rect 239 -160 241 -154
rect 249 -160 251 -154
rect 259 -160 261 -154
rect 291 -159 293 -145
rect 302 -165 304 -145
rect 309 -165 311 -145
rect 329 -165 331 -151
rect 339 -165 341 -151
rect 349 -158 351 -148
rect 359 -158 361 -145
rect 391 -159 393 -145
rect 402 -165 404 -145
rect 409 -165 411 -145
rect 429 -165 431 -151
rect 439 -165 441 -151
rect 449 -158 451 -148
rect 459 -158 461 -145
rect 483 -160 485 -154
rect 493 -160 495 -154
rect 503 -160 505 -154
rect 535 -159 537 -145
rect 546 -165 548 -145
rect 553 -165 555 -145
rect 573 -165 575 -151
rect 583 -165 585 -151
rect 593 -158 595 -148
rect 603 -158 605 -145
rect 635 -159 637 -145
rect 646 -165 648 -145
rect 653 -165 655 -145
rect 673 -165 675 -151
rect 683 -165 685 -151
rect 693 -158 695 -148
rect 703 -158 705 -145
rect 14 -277 16 -264
rect 24 -274 26 -264
rect 34 -271 36 -257
rect 44 -271 46 -257
rect 64 -277 66 -257
rect 71 -277 73 -257
rect 82 -277 84 -263
rect 114 -277 116 -264
rect 124 -274 126 -264
rect 134 -271 136 -257
rect 144 -271 146 -257
rect 164 -277 166 -257
rect 171 -277 173 -257
rect 182 -277 184 -263
rect 214 -268 216 -262
rect 224 -268 226 -262
rect 234 -268 236 -262
rect 255 -277 257 -264
rect 265 -274 267 -264
rect 275 -271 277 -257
rect 285 -271 287 -257
rect 305 -277 307 -257
rect 312 -277 314 -257
rect 323 -277 325 -263
rect 355 -277 357 -264
rect 365 -274 367 -264
rect 375 -271 377 -257
rect 385 -271 387 -257
rect 405 -277 407 -257
rect 412 -277 414 -257
rect 423 -277 425 -263
rect 455 -268 457 -262
rect 465 -268 467 -262
rect 475 -268 477 -262
<< pmos >>
rect 14 43 16 55
rect 24 43 26 53
rect 34 43 36 53
rect 58 43 60 55
rect 68 43 70 53
rect 78 43 80 53
rect 102 43 104 55
rect 112 43 114 53
rect 122 43 124 53
rect 146 43 148 55
rect 156 43 158 53
rect 166 43 168 53
rect 190 43 192 55
rect 200 43 202 53
rect 210 43 212 53
rect 234 43 236 55
rect 244 43 246 53
rect 254 43 256 53
rect 278 43 280 55
rect 288 43 290 53
rect 298 43 300 53
rect 322 43 324 55
rect 332 43 334 53
rect 342 43 344 53
rect 366 43 368 55
rect 376 43 378 53
rect 386 43 388 53
rect 410 43 412 55
rect 420 43 422 53
rect 430 43 432 53
rect 454 43 456 55
rect 464 43 466 53
rect 474 43 476 53
rect 498 43 500 55
rect 508 43 510 53
rect 518 43 520 53
rect 542 43 544 55
rect 552 43 554 53
rect 562 43 564 53
rect 586 43 588 55
rect 596 43 598 53
rect 606 43 608 53
rect 630 43 632 55
rect 640 43 642 53
rect 650 43 652 53
rect 674 43 676 55
rect 684 43 686 53
rect 694 43 696 53
rect 22 -61 24 -33
rect 32 -61 34 -33
rect 42 -61 44 -33
rect 60 -58 62 -33
rect 67 -58 69 -33
rect 77 -49 79 -36
rect 90 -61 92 -36
rect 111 -61 113 -33
rect 121 -61 123 -33
rect 131 -61 133 -33
rect 149 -58 151 -33
rect 156 -58 158 -33
rect 166 -49 168 -36
rect 179 -61 181 -36
rect 199 -61 201 -43
rect 206 -61 208 -43
rect 219 -52 221 -40
rect 240 -61 242 -33
rect 250 -61 252 -33
rect 260 -61 262 -33
rect 278 -58 280 -33
rect 285 -58 287 -33
rect 295 -49 297 -36
rect 308 -61 310 -36
rect 329 -61 331 -33
rect 339 -61 341 -33
rect 349 -61 351 -33
rect 367 -58 369 -33
rect 374 -58 376 -33
rect 384 -49 386 -36
rect 397 -61 399 -36
rect 498 -61 500 -33
rect 508 -61 510 -33
rect 518 -61 520 -33
rect 536 -58 538 -33
rect 543 -58 545 -33
rect 553 -49 555 -36
rect 566 -61 568 -36
rect 587 -61 589 -33
rect 597 -61 599 -33
rect 607 -61 609 -33
rect 625 -58 627 -33
rect 632 -58 634 -33
rect 642 -49 644 -36
rect 655 -61 657 -36
rect 14 -98 16 -73
rect 27 -98 29 -85
rect 37 -101 39 -76
rect 44 -101 46 -76
rect 62 -101 64 -73
rect 72 -101 74 -73
rect 82 -101 84 -73
rect 103 -98 105 -73
rect 116 -98 118 -85
rect 126 -101 128 -76
rect 133 -101 135 -76
rect 151 -101 153 -73
rect 161 -101 163 -73
rect 171 -101 173 -73
rect 192 -94 194 -82
rect 205 -91 207 -73
rect 212 -91 214 -73
rect 232 -98 234 -73
rect 245 -98 247 -85
rect 255 -101 257 -76
rect 262 -101 264 -76
rect 280 -101 282 -73
rect 290 -101 292 -73
rect 300 -101 302 -73
rect 321 -98 323 -73
rect 334 -98 336 -85
rect 344 -101 346 -76
rect 351 -101 353 -76
rect 369 -101 371 -73
rect 379 -101 381 -73
rect 389 -101 391 -73
rect 410 -94 412 -82
rect 423 -91 425 -73
rect 430 -91 432 -73
rect 450 -98 452 -73
rect 463 -98 465 -85
rect 473 -101 475 -76
rect 480 -101 482 -76
rect 498 -101 500 -73
rect 508 -101 510 -73
rect 518 -101 520 -73
rect 539 -98 541 -73
rect 552 -98 554 -85
rect 562 -101 564 -76
rect 569 -101 571 -76
rect 587 -101 589 -73
rect 597 -101 599 -73
rect 607 -101 609 -73
rect 628 -94 630 -82
rect 641 -91 643 -73
rect 648 -91 650 -73
rect 239 -205 241 -187
rect 246 -205 248 -187
rect 259 -196 261 -184
rect 291 -205 293 -177
rect 301 -205 303 -177
rect 311 -205 313 -177
rect 329 -202 331 -177
rect 336 -202 338 -177
rect 346 -193 348 -180
rect 359 -205 361 -180
rect 391 -205 393 -177
rect 401 -205 403 -177
rect 411 -205 413 -177
rect 429 -202 431 -177
rect 436 -202 438 -177
rect 446 -193 448 -180
rect 459 -205 461 -180
rect 483 -205 485 -187
rect 490 -205 492 -187
rect 503 -196 505 -184
rect 535 -205 537 -177
rect 545 -205 547 -177
rect 555 -205 557 -177
rect 573 -202 575 -177
rect 580 -202 582 -177
rect 590 -193 592 -180
rect 603 -205 605 -180
rect 635 -205 637 -177
rect 645 -205 647 -177
rect 655 -205 657 -177
rect 673 -202 675 -177
rect 680 -202 682 -177
rect 690 -193 692 -180
rect 703 -205 705 -180
rect 14 -242 16 -217
rect 27 -242 29 -229
rect 37 -245 39 -220
rect 44 -245 46 -220
rect 62 -245 64 -217
rect 72 -245 74 -217
rect 82 -245 84 -217
rect 114 -242 116 -217
rect 127 -242 129 -229
rect 137 -245 139 -220
rect 144 -245 146 -220
rect 162 -245 164 -217
rect 172 -245 174 -217
rect 182 -245 184 -217
rect 214 -238 216 -226
rect 227 -235 229 -217
rect 234 -235 236 -217
rect 255 -242 257 -217
rect 268 -242 270 -229
rect 278 -245 280 -220
rect 285 -245 287 -220
rect 303 -245 305 -217
rect 313 -245 315 -217
rect 323 -245 325 -217
rect 355 -242 357 -217
rect 368 -242 370 -229
rect 378 -245 380 -220
rect 385 -245 387 -220
rect 403 -245 405 -217
rect 413 -245 415 -217
rect 423 -245 425 -217
rect 455 -238 457 -226
rect 468 -235 470 -217
rect 475 -235 477 -217
<< polyct0 >>
rect 16 36 18 38
rect 60 36 62 38
rect 104 36 106 38
rect 148 36 150 38
rect 192 36 194 38
rect 236 36 238 38
rect 280 36 282 38
rect 324 36 326 38
rect 368 36 370 38
rect 412 36 414 38
rect 456 36 458 38
rect 500 36 502 38
rect 544 36 546 38
rect 588 36 590 38
rect 632 36 634 38
rect 676 36 678 38
rect 22 -28 24 -26
rect 32 -28 34 -26
rect 88 -21 90 -19
rect 82 -31 84 -29
rect 111 -28 113 -26
rect 121 -28 123 -26
rect 177 -21 179 -19
rect 171 -31 173 -29
rect 217 -29 219 -27
rect 240 -28 242 -26
rect 250 -28 252 -26
rect 306 -21 308 -19
rect 300 -31 302 -29
rect 329 -28 331 -26
rect 339 -28 341 -26
rect 395 -21 397 -19
rect 389 -31 391 -29
rect 498 -28 500 -26
rect 508 -28 510 -26
rect 564 -21 566 -19
rect 558 -31 560 -29
rect 587 -28 589 -26
rect 597 -28 599 -26
rect 653 -21 655 -19
rect 647 -31 649 -29
rect 22 -105 24 -103
rect 16 -115 18 -113
rect 72 -108 74 -106
rect 82 -108 84 -106
rect 111 -105 113 -103
rect 105 -115 107 -113
rect 161 -108 163 -106
rect 171 -108 173 -106
rect 194 -107 196 -105
rect 240 -105 242 -103
rect 234 -115 236 -113
rect 290 -108 292 -106
rect 300 -108 302 -106
rect 329 -105 331 -103
rect 323 -115 325 -113
rect 379 -108 381 -106
rect 389 -108 391 -106
rect 412 -107 414 -105
rect 458 -105 460 -103
rect 452 -115 454 -113
rect 508 -108 510 -106
rect 518 -108 520 -106
rect 547 -105 549 -103
rect 541 -115 543 -113
rect 597 -108 599 -106
rect 607 -108 609 -106
rect 630 -107 632 -105
rect 257 -173 259 -171
rect 291 -172 293 -170
rect 301 -172 303 -170
rect 357 -165 359 -163
rect 351 -175 353 -173
rect 391 -172 393 -170
rect 401 -172 403 -170
rect 457 -165 459 -163
rect 451 -175 453 -173
rect 501 -173 503 -171
rect 535 -172 537 -170
rect 545 -172 547 -170
rect 601 -165 603 -163
rect 595 -175 597 -173
rect 635 -172 637 -170
rect 645 -172 647 -170
rect 701 -165 703 -163
rect 695 -175 697 -173
rect 22 -249 24 -247
rect 16 -259 18 -257
rect 72 -252 74 -250
rect 82 -252 84 -250
rect 122 -249 124 -247
rect 116 -259 118 -257
rect 172 -252 174 -250
rect 182 -252 184 -250
rect 216 -251 218 -249
rect 263 -249 265 -247
rect 257 -259 259 -257
rect 313 -252 315 -250
rect 323 -252 325 -250
rect 363 -249 365 -247
rect 357 -259 359 -257
rect 413 -252 415 -250
rect 423 -252 425 -250
rect 457 -251 459 -249
<< polyct1 >>
rect 26 60 28 62
rect 70 60 72 62
rect 114 60 116 62
rect 158 60 160 62
rect 202 60 204 62
rect 246 60 248 62
rect 290 60 292 62
rect 334 60 336 62
rect 378 60 380 62
rect 422 60 424 62
rect 466 60 468 62
rect 510 60 512 62
rect 554 60 556 62
rect 598 60 600 62
rect 642 60 644 62
rect 686 60 688 62
rect 35 28 37 30
rect 79 28 81 30
rect 123 28 125 30
rect 167 28 169 30
rect 211 28 213 30
rect 255 28 257 30
rect 299 28 301 30
rect 343 28 345 30
rect 387 28 389 30
rect 431 28 433 30
rect 475 28 477 30
rect 519 28 521 30
rect 563 28 565 30
rect 607 28 609 30
rect 651 28 653 30
rect 695 28 697 30
rect 42 -28 44 -26
rect 49 -28 51 -26
rect 68 -28 70 -26
rect 131 -28 133 -26
rect 138 -28 140 -26
rect 157 -28 159 -26
rect 197 -28 199 -26
rect 260 -28 262 -26
rect 267 -28 269 -26
rect 286 -28 288 -26
rect 207 -36 209 -34
rect 349 -28 351 -26
rect 356 -28 358 -26
rect 375 -28 377 -26
rect 518 -28 520 -26
rect 525 -28 527 -26
rect 544 -28 546 -26
rect 607 -28 609 -26
rect 614 -28 616 -26
rect 633 -28 635 -26
rect 36 -108 38 -106
rect 55 -108 57 -106
rect 62 -108 64 -106
rect 204 -100 206 -98
rect 125 -108 127 -106
rect 144 -108 146 -106
rect 151 -108 153 -106
rect 214 -108 216 -106
rect 254 -108 256 -106
rect 273 -108 275 -106
rect 280 -108 282 -106
rect 422 -100 424 -98
rect 343 -108 345 -106
rect 362 -108 364 -106
rect 369 -108 371 -106
rect 432 -108 434 -106
rect 472 -108 474 -106
rect 491 -108 493 -106
rect 498 -108 500 -106
rect 640 -100 642 -98
rect 561 -108 563 -106
rect 580 -108 582 -106
rect 587 -108 589 -106
rect 650 -108 652 -106
rect 237 -172 239 -170
rect 311 -172 313 -170
rect 318 -172 320 -170
rect 337 -172 339 -170
rect 247 -180 249 -178
rect 411 -172 413 -170
rect 418 -172 420 -170
rect 437 -172 439 -170
rect 481 -172 483 -170
rect 555 -172 557 -170
rect 562 -172 564 -170
rect 581 -172 583 -170
rect 491 -180 493 -178
rect 655 -172 657 -170
rect 662 -172 664 -170
rect 681 -172 683 -170
rect 36 -252 38 -250
rect 55 -252 57 -250
rect 62 -252 64 -250
rect 226 -244 228 -242
rect 136 -252 138 -250
rect 155 -252 157 -250
rect 162 -252 164 -250
rect 236 -252 238 -250
rect 277 -252 279 -250
rect 296 -252 298 -250
rect 303 -252 305 -250
rect 467 -244 469 -242
rect 377 -252 379 -250
rect 396 -252 398 -250
rect 403 -252 405 -250
rect 477 -252 479 -250
<< ndifct0 >>
rect 38 19 40 21
rect 82 19 84 21
rect 126 19 128 21
rect 170 19 172 21
rect 214 19 216 21
rect 258 19 260 21
rect 302 19 304 21
rect 346 19 348 21
rect 390 19 392 21
rect 434 19 436 21
rect 478 19 480 21
rect 522 19 524 21
rect 566 19 568 21
rect 610 19 612 21
rect 654 19 656 21
rect 698 19 700 21
rect 28 -5 30 -3
rect 45 -12 47 -10
rect 55 -12 57 -10
rect 55 -19 57 -17
rect 65 -19 67 -17
rect 75 -11 77 -9
rect 85 -8 87 -6
rect 117 -5 119 -3
rect 134 -12 136 -10
rect 144 -12 146 -10
rect 144 -19 146 -17
rect 154 -19 156 -17
rect 164 -11 166 -9
rect 174 -8 176 -6
rect 194 -14 196 -12
rect 204 -14 206 -12
rect 214 -14 216 -12
rect 246 -5 248 -3
rect 263 -12 265 -10
rect 273 -12 275 -10
rect 273 -19 275 -17
rect 283 -19 285 -17
rect 293 -11 295 -9
rect 303 -8 305 -6
rect 335 -5 337 -3
rect 352 -12 354 -10
rect 362 -12 364 -10
rect 362 -19 364 -17
rect 372 -19 374 -17
rect 382 -11 384 -9
rect 392 -8 394 -6
rect 504 -5 506 -3
rect 521 -12 523 -10
rect 531 -12 533 -10
rect 531 -19 533 -17
rect 541 -19 543 -17
rect 551 -11 553 -9
rect 561 -8 563 -6
rect 593 -5 595 -3
rect 610 -12 612 -10
rect 620 -12 622 -10
rect 620 -19 622 -17
rect 630 -19 632 -17
rect 640 -11 642 -9
rect 650 -8 652 -6
rect 19 -128 21 -126
rect 29 -125 31 -123
rect 39 -117 41 -115
rect 49 -117 51 -115
rect 49 -124 51 -122
rect 59 -124 61 -122
rect 76 -131 78 -129
rect 108 -128 110 -126
rect 118 -125 120 -123
rect 128 -117 130 -115
rect 138 -117 140 -115
rect 138 -124 140 -122
rect 148 -124 150 -122
rect 165 -131 167 -129
rect 197 -122 199 -120
rect 207 -122 209 -120
rect 217 -122 219 -120
rect 237 -128 239 -126
rect 247 -125 249 -123
rect 257 -117 259 -115
rect 267 -117 269 -115
rect 267 -124 269 -122
rect 277 -124 279 -122
rect 294 -131 296 -129
rect 326 -128 328 -126
rect 336 -125 338 -123
rect 346 -117 348 -115
rect 356 -117 358 -115
rect 356 -124 358 -122
rect 366 -124 368 -122
rect 383 -131 385 -129
rect 415 -122 417 -120
rect 425 -122 427 -120
rect 435 -122 437 -120
rect 455 -128 457 -126
rect 465 -125 467 -123
rect 475 -117 477 -115
rect 485 -117 487 -115
rect 485 -124 487 -122
rect 495 -124 497 -122
rect 512 -131 514 -129
rect 544 -128 546 -126
rect 554 -125 556 -123
rect 564 -117 566 -115
rect 574 -117 576 -115
rect 574 -124 576 -122
rect 584 -124 586 -122
rect 601 -131 603 -129
rect 633 -122 635 -120
rect 643 -122 645 -120
rect 653 -122 655 -120
rect 234 -158 236 -156
rect 244 -158 246 -156
rect 254 -158 256 -156
rect 297 -149 299 -147
rect 314 -156 316 -154
rect 324 -156 326 -154
rect 324 -163 326 -161
rect 334 -163 336 -161
rect 344 -155 346 -153
rect 354 -152 356 -150
rect 397 -149 399 -147
rect 414 -156 416 -154
rect 424 -156 426 -154
rect 424 -163 426 -161
rect 434 -163 436 -161
rect 444 -155 446 -153
rect 454 -152 456 -150
rect 478 -158 480 -156
rect 488 -158 490 -156
rect 498 -158 500 -156
rect 541 -149 543 -147
rect 558 -156 560 -154
rect 568 -156 570 -154
rect 568 -163 570 -161
rect 578 -163 580 -161
rect 588 -155 590 -153
rect 598 -152 600 -150
rect 641 -149 643 -147
rect 658 -156 660 -154
rect 668 -156 670 -154
rect 668 -163 670 -161
rect 678 -163 680 -161
rect 688 -155 690 -153
rect 698 -152 700 -150
rect 19 -272 21 -270
rect 29 -269 31 -267
rect 39 -261 41 -259
rect 49 -261 51 -259
rect 49 -268 51 -266
rect 59 -268 61 -266
rect 76 -275 78 -273
rect 119 -272 121 -270
rect 129 -269 131 -267
rect 139 -261 141 -259
rect 149 -261 151 -259
rect 149 -268 151 -266
rect 159 -268 161 -266
rect 176 -275 178 -273
rect 219 -266 221 -264
rect 229 -266 231 -264
rect 239 -266 241 -264
rect 260 -272 262 -270
rect 270 -269 272 -267
rect 280 -261 282 -259
rect 290 -261 292 -259
rect 290 -268 292 -266
rect 300 -268 302 -266
rect 317 -275 319 -273
rect 360 -272 362 -270
rect 370 -269 372 -267
rect 380 -261 382 -259
rect 390 -261 392 -259
rect 390 -268 392 -266
rect 400 -268 402 -266
rect 417 -275 419 -273
rect 460 -266 462 -264
rect 470 -266 472 -264
rect 480 -266 482 -264
<< ndifct1 >>
rect 9 22 11 24
rect 53 22 55 24
rect 97 22 99 24
rect 141 22 143 24
rect 185 22 187 24
rect 229 22 231 24
rect 273 22 275 24
rect 317 22 319 24
rect 361 22 363 24
rect 405 22 407 24
rect 449 22 451 24
rect 493 22 495 24
rect 537 22 539 24
rect 581 22 583 24
rect 625 22 627 24
rect 669 22 671 24
rect 20 10 22 12
rect 64 10 66 12
rect 108 10 110 12
rect 152 10 154 12
rect 196 10 198 12
rect 240 10 242 12
rect 284 10 286 12
rect 328 10 330 12
rect 372 10 374 12
rect 416 10 418 12
rect 460 10 462 12
rect 504 10 506 12
rect 548 10 550 12
rect 592 10 594 12
rect 636 10 638 12
rect 680 10 682 12
rect 17 -12 19 -10
rect 95 -12 97 -10
rect 106 -12 108 -10
rect 184 -12 186 -10
rect 224 -14 226 -12
rect 235 -12 237 -10
rect 313 -12 315 -10
rect 324 -12 326 -10
rect 402 -12 404 -10
rect 493 -12 495 -10
rect 571 -12 573 -10
rect 582 -12 584 -10
rect 660 -12 662 -10
rect 9 -124 11 -122
rect 87 -124 89 -122
rect 98 -124 100 -122
rect 176 -124 178 -122
rect 187 -122 189 -120
rect 227 -124 229 -122
rect 305 -124 307 -122
rect 316 -124 318 -122
rect 394 -124 396 -122
rect 405 -122 407 -120
rect 445 -124 447 -122
rect 523 -124 525 -122
rect 534 -124 536 -122
rect 612 -124 614 -122
rect 623 -122 625 -120
rect 264 -158 266 -156
rect 286 -156 288 -154
rect 364 -156 366 -154
rect 386 -156 388 -154
rect 464 -156 466 -154
rect 508 -158 510 -156
rect 530 -156 532 -154
rect 608 -156 610 -154
rect 630 -156 632 -154
rect 708 -156 710 -154
rect 9 -268 11 -266
rect 87 -268 89 -266
rect 109 -268 111 -266
rect 187 -268 189 -266
rect 209 -266 211 -264
rect 250 -268 252 -266
rect 328 -268 330 -266
rect 350 -268 352 -266
rect 428 -268 430 -266
rect 450 -266 452 -264
<< ntiect1 >>
rect 10 70 12 72
rect 24 70 26 72
rect 38 70 40 72
rect 54 70 56 72
rect 68 70 70 72
rect 82 70 84 72
rect 98 70 100 72
rect 112 70 114 72
rect 126 70 128 72
rect 142 70 144 72
rect 156 70 158 72
rect 170 70 172 72
rect 186 70 188 72
rect 200 70 202 72
rect 214 70 216 72
rect 230 70 232 72
rect 244 70 246 72
rect 258 70 260 72
rect 274 70 276 72
rect 288 70 290 72
rect 302 70 304 72
rect 318 70 320 72
rect 332 70 334 72
rect 346 70 348 72
rect 362 70 364 72
rect 376 70 378 72
rect 390 70 392 72
rect 406 70 408 72
rect 420 70 422 72
rect 434 70 436 72
rect 450 70 452 72
rect 464 70 466 72
rect 478 70 480 72
rect 494 70 496 72
rect 508 70 510 72
rect 522 70 524 72
rect 538 70 540 72
rect 552 70 554 72
rect 566 70 568 72
rect 582 70 584 72
rect 596 70 598 72
rect 610 70 612 72
rect 626 70 628 72
rect 640 70 642 72
rect 654 70 656 72
rect 670 70 672 72
rect 684 70 686 72
rect 698 70 700 72
rect 223 -62 225 -60
rect 188 -74 190 -72
rect 406 -74 408 -72
rect 624 -74 626 -72
rect 263 -206 265 -204
rect 507 -206 509 -204
rect 210 -218 212 -216
rect 451 -218 453 -216
<< ptiect1 >>
rect 10 10 12 12
rect 54 10 56 12
rect 98 10 100 12
rect 142 10 144 12
rect 186 10 188 12
rect 230 10 232 12
rect 274 10 276 12
rect 318 10 320 12
rect 362 10 364 12
rect 406 10 408 12
rect 450 10 452 12
rect 494 10 496 12
rect 538 10 540 12
rect 582 10 584 12
rect 626 10 628 12
rect 670 10 672 12
rect 195 -2 197 0
rect 223 -2 225 0
rect 188 -134 190 -132
rect 216 -134 218 -132
rect 406 -134 408 -132
rect 434 -134 436 -132
rect 624 -134 626 -132
rect 652 -134 654 -132
rect 235 -146 237 -144
rect 263 -146 265 -144
rect 479 -146 481 -144
rect 507 -146 509 -144
rect 210 -278 212 -276
rect 238 -278 240 -276
rect 451 -278 453 -276
rect 479 -278 481 -276
<< pdifct0 >>
rect 19 45 21 47
rect 29 45 31 47
rect 39 49 41 51
rect 63 45 65 47
rect 73 45 75 47
rect 83 49 85 51
rect 107 45 109 47
rect 117 45 119 47
rect 127 49 129 51
rect 151 45 153 47
rect 161 45 163 47
rect 171 49 173 51
rect 195 45 197 47
rect 205 45 207 47
rect 215 49 217 51
rect 239 45 241 47
rect 249 45 251 47
rect 259 49 261 51
rect 283 45 285 47
rect 293 45 295 47
rect 303 49 305 51
rect 327 45 329 47
rect 337 45 339 47
rect 347 49 349 51
rect 371 45 373 47
rect 381 45 383 47
rect 391 49 393 51
rect 415 45 417 47
rect 425 45 427 47
rect 435 49 437 51
rect 459 45 461 47
rect 469 45 471 47
rect 479 49 481 51
rect 503 45 505 47
rect 513 45 515 47
rect 523 49 525 51
rect 547 45 549 47
rect 557 45 559 47
rect 567 49 569 51
rect 591 45 593 47
rect 601 45 603 47
rect 611 49 613 51
rect 635 45 637 47
rect 645 45 647 47
rect 655 49 657 51
rect 679 45 681 47
rect 689 45 691 47
rect 699 49 701 51
rect 27 -52 29 -50
rect 27 -59 29 -57
rect 37 -44 39 -42
rect 37 -51 39 -49
rect 49 -52 51 -50
rect 49 -59 51 -57
rect 72 -40 74 -38
rect 84 -59 86 -57
rect 116 -52 118 -50
rect 116 -59 118 -57
rect 126 -44 128 -42
rect 126 -51 128 -49
rect 138 -52 140 -50
rect 138 -59 140 -57
rect 161 -40 163 -38
rect 173 -59 175 -57
rect 194 -52 196 -50
rect 212 -59 214 -57
rect 245 -52 247 -50
rect 245 -59 247 -57
rect 255 -44 257 -42
rect 255 -51 257 -49
rect 267 -52 269 -50
rect 267 -59 269 -57
rect 290 -40 292 -38
rect 302 -59 304 -57
rect 334 -52 336 -50
rect 334 -59 336 -57
rect 344 -44 346 -42
rect 344 -51 346 -49
rect 356 -52 358 -50
rect 356 -59 358 -57
rect 379 -40 381 -38
rect 391 -59 393 -57
rect 503 -52 505 -50
rect 503 -59 505 -57
rect 513 -44 515 -42
rect 513 -51 515 -49
rect 525 -52 527 -50
rect 525 -59 527 -57
rect 548 -40 550 -38
rect 560 -59 562 -57
rect 592 -52 594 -50
rect 592 -59 594 -57
rect 602 -44 604 -42
rect 602 -51 604 -49
rect 614 -52 616 -50
rect 614 -59 616 -57
rect 637 -40 639 -38
rect 649 -59 651 -57
rect 20 -77 22 -75
rect 32 -96 34 -94
rect 55 -77 57 -75
rect 55 -84 57 -82
rect 67 -85 69 -83
rect 67 -92 69 -90
rect 77 -77 79 -75
rect 77 -84 79 -82
rect 109 -77 111 -75
rect 121 -96 123 -94
rect 144 -77 146 -75
rect 144 -84 146 -82
rect 156 -85 158 -83
rect 156 -92 158 -90
rect 166 -77 168 -75
rect 166 -84 168 -82
rect 199 -77 201 -75
rect 217 -84 219 -82
rect 238 -77 240 -75
rect 250 -96 252 -94
rect 273 -77 275 -75
rect 273 -84 275 -82
rect 285 -85 287 -83
rect 285 -92 287 -90
rect 295 -77 297 -75
rect 295 -84 297 -82
rect 327 -77 329 -75
rect 339 -96 341 -94
rect 362 -77 364 -75
rect 362 -84 364 -82
rect 374 -85 376 -83
rect 374 -92 376 -90
rect 384 -77 386 -75
rect 384 -84 386 -82
rect 417 -77 419 -75
rect 435 -84 437 -82
rect 456 -77 458 -75
rect 468 -96 470 -94
rect 491 -77 493 -75
rect 491 -84 493 -82
rect 503 -85 505 -83
rect 503 -92 505 -90
rect 513 -77 515 -75
rect 513 -84 515 -82
rect 545 -77 547 -75
rect 557 -96 559 -94
rect 580 -77 582 -75
rect 580 -84 582 -82
rect 592 -85 594 -83
rect 592 -92 594 -90
rect 602 -77 604 -75
rect 602 -84 604 -82
rect 635 -77 637 -75
rect 653 -84 655 -82
rect 234 -196 236 -194
rect 252 -203 254 -201
rect 296 -196 298 -194
rect 296 -203 298 -201
rect 306 -188 308 -186
rect 306 -195 308 -193
rect 318 -196 320 -194
rect 318 -203 320 -201
rect 341 -184 343 -182
rect 353 -203 355 -201
rect 396 -196 398 -194
rect 396 -203 398 -201
rect 406 -188 408 -186
rect 406 -195 408 -193
rect 418 -196 420 -194
rect 418 -203 420 -201
rect 441 -184 443 -182
rect 453 -203 455 -201
rect 478 -196 480 -194
rect 496 -203 498 -201
rect 540 -196 542 -194
rect 540 -203 542 -201
rect 550 -188 552 -186
rect 550 -195 552 -193
rect 562 -196 564 -194
rect 562 -203 564 -201
rect 585 -184 587 -182
rect 597 -203 599 -201
rect 640 -196 642 -194
rect 640 -203 642 -201
rect 650 -188 652 -186
rect 650 -195 652 -193
rect 662 -196 664 -194
rect 662 -203 664 -201
rect 685 -184 687 -182
rect 697 -203 699 -201
rect 20 -221 22 -219
rect 32 -240 34 -238
rect 55 -221 57 -219
rect 55 -228 57 -226
rect 67 -229 69 -227
rect 67 -236 69 -234
rect 77 -221 79 -219
rect 77 -228 79 -226
rect 120 -221 122 -219
rect 132 -240 134 -238
rect 155 -221 157 -219
rect 155 -228 157 -226
rect 167 -229 169 -227
rect 167 -236 169 -234
rect 177 -221 179 -219
rect 177 -228 179 -226
rect 221 -221 223 -219
rect 239 -228 241 -226
rect 261 -221 263 -219
rect 273 -240 275 -238
rect 296 -221 298 -219
rect 296 -228 298 -226
rect 308 -229 310 -227
rect 308 -236 310 -234
rect 318 -221 320 -219
rect 318 -228 320 -226
rect 361 -221 363 -219
rect 373 -240 375 -238
rect 396 -221 398 -219
rect 396 -228 398 -226
rect 408 -229 410 -227
rect 408 -236 410 -234
rect 418 -221 420 -219
rect 418 -228 420 -226
rect 462 -221 464 -219
rect 480 -228 482 -226
<< pdifct1 >>
rect 9 45 11 47
rect 53 45 55 47
rect 97 45 99 47
rect 141 45 143 47
rect 185 45 187 47
rect 229 45 231 47
rect 273 45 275 47
rect 317 45 319 47
rect 361 45 363 47
rect 405 45 407 47
rect 449 45 451 47
rect 493 45 495 47
rect 537 45 539 47
rect 581 45 583 47
rect 625 45 627 47
rect 669 45 671 47
rect 17 -37 19 -35
rect 17 -44 19 -42
rect 95 -40 97 -38
rect 95 -47 97 -45
rect 106 -37 108 -35
rect 106 -44 108 -42
rect 184 -40 186 -38
rect 235 -37 237 -35
rect 184 -47 186 -45
rect 235 -44 237 -42
rect 224 -50 226 -48
rect 313 -40 315 -38
rect 313 -47 315 -45
rect 324 -37 326 -35
rect 324 -44 326 -42
rect 402 -40 404 -38
rect 402 -47 404 -45
rect 493 -37 495 -35
rect 493 -44 495 -42
rect 571 -40 573 -38
rect 571 -47 573 -45
rect 582 -37 584 -35
rect 582 -44 584 -42
rect 660 -40 662 -38
rect 660 -47 662 -45
rect 9 -89 11 -87
rect 9 -96 11 -94
rect 87 -92 89 -90
rect 87 -99 89 -97
rect 98 -89 100 -87
rect 98 -96 100 -94
rect 187 -86 189 -84
rect 176 -92 178 -90
rect 227 -89 229 -87
rect 176 -99 178 -97
rect 227 -96 229 -94
rect 305 -92 307 -90
rect 305 -99 307 -97
rect 316 -89 318 -87
rect 316 -96 318 -94
rect 405 -86 407 -84
rect 394 -92 396 -90
rect 445 -89 447 -87
rect 394 -99 396 -97
rect 445 -96 447 -94
rect 523 -92 525 -90
rect 523 -99 525 -97
rect 534 -89 536 -87
rect 534 -96 536 -94
rect 623 -86 625 -84
rect 612 -92 614 -90
rect 612 -99 614 -97
rect 286 -181 288 -179
rect 286 -188 288 -186
rect 264 -194 266 -192
rect 364 -184 366 -182
rect 364 -191 366 -189
rect 386 -181 388 -179
rect 386 -188 388 -186
rect 464 -184 466 -182
rect 530 -181 532 -179
rect 464 -191 466 -189
rect 530 -188 532 -186
rect 508 -194 510 -192
rect 608 -184 610 -182
rect 608 -191 610 -189
rect 630 -181 632 -179
rect 630 -188 632 -186
rect 708 -184 710 -182
rect 708 -191 710 -189
rect 9 -233 11 -231
rect 9 -240 11 -238
rect 87 -236 89 -234
rect 87 -243 89 -241
rect 109 -233 111 -231
rect 109 -240 111 -238
rect 209 -230 211 -228
rect 187 -236 189 -234
rect 250 -233 252 -231
rect 187 -243 189 -241
rect 250 -240 252 -238
rect 328 -236 330 -234
rect 328 -243 330 -241
rect 350 -233 352 -231
rect 350 -240 352 -238
rect 450 -230 452 -228
rect 428 -236 430 -234
rect 428 -243 430 -241
<< alu0 >>
rect 11 43 12 49
rect 15 48 19 69
rect 38 51 42 69
rect 38 49 39 51
rect 41 49 42 51
rect 15 47 23 48
rect 15 45 19 47
rect 21 45 23 47
rect 15 44 23 45
rect 27 47 33 48
rect 38 47 42 49
rect 27 45 29 47
rect 31 45 33 47
rect 27 39 33 45
rect 14 38 33 39
rect 14 36 16 38
rect 18 36 33 38
rect 14 35 33 36
rect 11 24 12 26
rect 23 22 27 35
rect 55 43 56 49
rect 59 48 63 69
rect 82 51 86 69
rect 82 49 83 51
rect 85 49 86 51
rect 59 47 67 48
rect 59 45 63 47
rect 65 45 67 47
rect 59 44 67 45
rect 71 47 77 48
rect 82 47 86 49
rect 71 45 73 47
rect 75 45 77 47
rect 71 39 77 45
rect 58 38 77 39
rect 58 36 60 38
rect 62 36 77 38
rect 58 35 77 36
rect 55 24 56 26
rect 23 21 42 22
rect 23 19 38 21
rect 40 19 42 21
rect 23 18 42 19
rect 67 22 71 35
rect 99 43 100 49
rect 103 48 107 69
rect 126 51 130 69
rect 126 49 127 51
rect 129 49 130 51
rect 103 47 111 48
rect 103 45 107 47
rect 109 45 111 47
rect 103 44 111 45
rect 115 47 121 48
rect 126 47 130 49
rect 115 45 117 47
rect 119 45 121 47
rect 115 39 121 45
rect 102 38 121 39
rect 102 36 104 38
rect 106 36 121 38
rect 102 35 121 36
rect 99 24 100 26
rect 67 21 86 22
rect 67 19 82 21
rect 84 19 86 21
rect 67 18 86 19
rect 111 22 115 35
rect 143 43 144 49
rect 147 48 151 69
rect 170 51 174 69
rect 170 49 171 51
rect 173 49 174 51
rect 147 47 155 48
rect 147 45 151 47
rect 153 45 155 47
rect 147 44 155 45
rect 159 47 165 48
rect 170 47 174 49
rect 159 45 161 47
rect 163 45 165 47
rect 159 39 165 45
rect 146 38 165 39
rect 146 36 148 38
rect 150 36 165 38
rect 146 35 165 36
rect 143 24 144 26
rect 111 21 130 22
rect 111 19 126 21
rect 128 19 130 21
rect 111 18 130 19
rect 155 22 159 35
rect 187 43 188 49
rect 191 48 195 69
rect 214 51 218 69
rect 214 49 215 51
rect 217 49 218 51
rect 191 47 199 48
rect 191 45 195 47
rect 197 45 199 47
rect 191 44 199 45
rect 203 47 209 48
rect 214 47 218 49
rect 203 45 205 47
rect 207 45 209 47
rect 203 39 209 45
rect 190 38 209 39
rect 190 36 192 38
rect 194 36 209 38
rect 190 35 209 36
rect 187 24 188 26
rect 155 21 174 22
rect 155 19 170 21
rect 172 19 174 21
rect 155 18 174 19
rect 199 22 203 35
rect 231 43 232 49
rect 235 48 239 69
rect 258 51 262 69
rect 258 49 259 51
rect 261 49 262 51
rect 235 47 243 48
rect 235 45 239 47
rect 241 45 243 47
rect 235 44 243 45
rect 247 47 253 48
rect 258 47 262 49
rect 247 45 249 47
rect 251 45 253 47
rect 247 39 253 45
rect 234 38 253 39
rect 234 36 236 38
rect 238 36 253 38
rect 234 35 253 36
rect 231 24 232 26
rect 199 21 218 22
rect 199 19 214 21
rect 216 19 218 21
rect 199 18 218 19
rect 243 22 247 35
rect 275 43 276 49
rect 279 48 283 69
rect 302 51 306 69
rect 302 49 303 51
rect 305 49 306 51
rect 279 47 287 48
rect 279 45 283 47
rect 285 45 287 47
rect 279 44 287 45
rect 291 47 297 48
rect 302 47 306 49
rect 291 45 293 47
rect 295 45 297 47
rect 291 39 297 45
rect 278 38 297 39
rect 278 36 280 38
rect 282 36 297 38
rect 278 35 297 36
rect 275 24 276 26
rect 243 21 262 22
rect 243 19 258 21
rect 260 19 262 21
rect 243 18 262 19
rect 287 22 291 35
rect 319 43 320 49
rect 323 48 327 69
rect 346 51 350 69
rect 346 49 347 51
rect 349 49 350 51
rect 323 47 331 48
rect 323 45 327 47
rect 329 45 331 47
rect 323 44 331 45
rect 335 47 341 48
rect 346 47 350 49
rect 335 45 337 47
rect 339 45 341 47
rect 335 39 341 45
rect 322 38 341 39
rect 322 36 324 38
rect 326 36 341 38
rect 322 35 341 36
rect 319 24 320 26
rect 287 21 306 22
rect 287 19 302 21
rect 304 19 306 21
rect 287 18 306 19
rect 331 22 335 35
rect 363 43 364 49
rect 367 48 371 69
rect 390 51 394 69
rect 390 49 391 51
rect 393 49 394 51
rect 367 47 375 48
rect 367 45 371 47
rect 373 45 375 47
rect 367 44 375 45
rect 379 47 385 48
rect 390 47 394 49
rect 379 45 381 47
rect 383 45 385 47
rect 379 39 385 45
rect 366 38 385 39
rect 366 36 368 38
rect 370 36 385 38
rect 366 35 385 36
rect 363 24 364 26
rect 331 21 350 22
rect 331 19 346 21
rect 348 19 350 21
rect 331 18 350 19
rect 375 22 379 35
rect 407 43 408 49
rect 411 48 415 69
rect 434 51 438 69
rect 434 49 435 51
rect 437 49 438 51
rect 411 47 419 48
rect 411 45 415 47
rect 417 45 419 47
rect 411 44 419 45
rect 423 47 429 48
rect 434 47 438 49
rect 423 45 425 47
rect 427 45 429 47
rect 423 39 429 45
rect 410 38 429 39
rect 410 36 412 38
rect 414 36 429 38
rect 410 35 429 36
rect 407 24 408 26
rect 375 21 394 22
rect 375 19 390 21
rect 392 19 394 21
rect 375 18 394 19
rect 419 22 423 35
rect 451 43 452 49
rect 455 48 459 69
rect 478 51 482 69
rect 478 49 479 51
rect 481 49 482 51
rect 455 47 463 48
rect 455 45 459 47
rect 461 45 463 47
rect 455 44 463 45
rect 467 47 473 48
rect 478 47 482 49
rect 467 45 469 47
rect 471 45 473 47
rect 467 39 473 45
rect 454 38 473 39
rect 454 36 456 38
rect 458 36 473 38
rect 454 35 473 36
rect 451 24 452 26
rect 419 21 438 22
rect 419 19 434 21
rect 436 19 438 21
rect 419 18 438 19
rect 463 22 467 35
rect 495 43 496 49
rect 499 48 503 69
rect 522 51 526 69
rect 522 49 523 51
rect 525 49 526 51
rect 499 47 507 48
rect 499 45 503 47
rect 505 45 507 47
rect 499 44 507 45
rect 511 47 517 48
rect 522 47 526 49
rect 511 45 513 47
rect 515 45 517 47
rect 511 39 517 45
rect 498 38 517 39
rect 498 36 500 38
rect 502 36 517 38
rect 498 35 517 36
rect 495 24 496 26
rect 463 21 482 22
rect 463 19 478 21
rect 480 19 482 21
rect 463 18 482 19
rect 507 22 511 35
rect 539 43 540 49
rect 543 48 547 69
rect 566 51 570 69
rect 566 49 567 51
rect 569 49 570 51
rect 543 47 551 48
rect 543 45 547 47
rect 549 45 551 47
rect 543 44 551 45
rect 555 47 561 48
rect 566 47 570 49
rect 555 45 557 47
rect 559 45 561 47
rect 555 39 561 45
rect 542 38 561 39
rect 542 36 544 38
rect 546 36 561 38
rect 542 35 561 36
rect 539 24 540 26
rect 507 21 526 22
rect 507 19 522 21
rect 524 19 526 21
rect 507 18 526 19
rect 551 22 555 35
rect 583 43 584 49
rect 587 48 591 69
rect 610 51 614 69
rect 610 49 611 51
rect 613 49 614 51
rect 587 47 595 48
rect 587 45 591 47
rect 593 45 595 47
rect 587 44 595 45
rect 599 47 605 48
rect 610 47 614 49
rect 599 45 601 47
rect 603 45 605 47
rect 599 39 605 45
rect 586 38 605 39
rect 586 36 588 38
rect 590 36 605 38
rect 586 35 605 36
rect 583 24 584 26
rect 551 21 570 22
rect 551 19 566 21
rect 568 19 570 21
rect 551 18 570 19
rect 595 22 599 35
rect 627 43 628 49
rect 631 48 635 69
rect 654 51 658 69
rect 654 49 655 51
rect 657 49 658 51
rect 631 47 639 48
rect 631 45 635 47
rect 637 45 639 47
rect 631 44 639 45
rect 643 47 649 48
rect 654 47 658 49
rect 643 45 645 47
rect 647 45 649 47
rect 643 39 649 45
rect 630 38 649 39
rect 630 36 632 38
rect 634 36 649 38
rect 630 35 649 36
rect 627 24 628 26
rect 595 21 614 22
rect 595 19 610 21
rect 612 19 614 21
rect 595 18 614 19
rect 639 22 643 35
rect 671 43 672 49
rect 675 48 679 69
rect 698 51 702 69
rect 698 49 699 51
rect 701 49 702 51
rect 675 47 683 48
rect 675 45 679 47
rect 681 45 683 47
rect 675 44 683 45
rect 687 47 693 48
rect 698 47 702 49
rect 687 45 689 47
rect 691 45 693 47
rect 687 39 693 45
rect 674 38 693 39
rect 674 36 676 38
rect 678 36 693 38
rect 674 35 693 36
rect 671 24 672 26
rect 639 21 658 22
rect 639 19 654 21
rect 656 19 658 21
rect 639 18 658 19
rect 683 22 687 35
rect 683 21 702 22
rect 683 19 698 21
rect 700 19 702 21
rect 683 18 702 19
rect 26 -5 28 -3
rect 30 -5 32 -3
rect 26 -6 32 -5
rect 84 -6 88 -3
rect 115 -5 117 -3
rect 119 -5 121 -3
rect 115 -6 121 -5
rect 173 -6 177 -3
rect 84 -8 85 -6
rect 87 -8 88 -6
rect 173 -8 174 -6
rect 176 -8 177 -6
rect 54 -9 79 -8
rect 39 -10 49 -9
rect 39 -12 45 -10
rect 47 -12 49 -10
rect 39 -13 49 -12
rect 54 -10 75 -9
rect 54 -12 55 -10
rect 57 -11 75 -10
rect 77 -11 79 -9
rect 84 -10 88 -8
rect 143 -9 168 -8
rect 57 -12 79 -11
rect 39 -17 43 -13
rect 23 -21 43 -17
rect 23 -24 27 -21
rect 21 -26 27 -24
rect 21 -28 22 -26
rect 24 -28 27 -26
rect 21 -30 27 -28
rect 23 -41 27 -30
rect 31 -26 35 -24
rect 54 -17 58 -12
rect 54 -19 55 -17
rect 57 -19 58 -17
rect 54 -21 58 -19
rect 63 -17 78 -16
rect 63 -19 65 -17
rect 67 -18 78 -17
rect 67 -19 92 -18
rect 63 -20 88 -19
rect 74 -21 88 -20
rect 90 -21 92 -19
rect 74 -22 92 -21
rect 31 -28 32 -26
rect 34 -28 35 -26
rect 31 -33 35 -28
rect 74 -33 78 -22
rect 71 -37 78 -33
rect 81 -29 85 -27
rect 81 -31 82 -29
rect 84 -31 85 -29
rect 71 -38 75 -37
rect 71 -40 72 -38
rect 74 -40 75 -38
rect 23 -42 63 -41
rect 71 -42 75 -40
rect 81 -41 85 -31
rect 23 -44 37 -42
rect 39 -44 63 -42
rect 23 -45 63 -44
rect 79 -45 85 -41
rect 36 -49 40 -45
rect 59 -49 83 -45
rect 128 -10 138 -9
rect 128 -12 134 -10
rect 136 -12 138 -10
rect 128 -13 138 -12
rect 143 -10 164 -9
rect 143 -12 144 -10
rect 146 -11 164 -10
rect 166 -11 168 -9
rect 173 -10 177 -8
rect 146 -12 168 -11
rect 128 -17 132 -13
rect 112 -21 132 -17
rect 112 -24 116 -21
rect 110 -26 116 -24
rect 110 -28 111 -26
rect 113 -28 116 -26
rect 110 -30 116 -28
rect 112 -41 116 -30
rect 120 -26 124 -24
rect 143 -17 147 -12
rect 143 -19 144 -17
rect 146 -19 147 -17
rect 143 -21 147 -19
rect 152 -17 167 -16
rect 152 -19 154 -17
rect 156 -18 167 -17
rect 192 -12 198 -3
rect 192 -14 194 -12
rect 196 -14 198 -12
rect 192 -15 198 -14
rect 203 -12 207 -10
rect 203 -14 204 -12
rect 206 -14 207 -12
rect 156 -19 181 -18
rect 152 -20 177 -19
rect 163 -21 177 -20
rect 179 -21 181 -19
rect 163 -22 181 -21
rect 120 -28 121 -26
rect 123 -28 124 -26
rect 120 -33 124 -28
rect 163 -33 167 -22
rect 160 -37 167 -33
rect 170 -29 174 -27
rect 170 -31 171 -29
rect 173 -31 174 -29
rect 160 -38 164 -37
rect 160 -40 161 -38
rect 163 -40 164 -38
rect 112 -42 152 -41
rect 160 -42 164 -40
rect 170 -41 174 -31
rect 203 -18 207 -14
rect 212 -12 218 -3
rect 244 -5 246 -3
rect 248 -5 250 -3
rect 244 -6 250 -5
rect 302 -6 306 -3
rect 333 -5 335 -3
rect 337 -5 339 -3
rect 333 -6 339 -5
rect 391 -6 395 -3
rect 502 -5 504 -3
rect 506 -5 508 -3
rect 502 -6 508 -5
rect 560 -6 564 -3
rect 591 -5 593 -3
rect 595 -5 597 -3
rect 591 -6 597 -5
rect 649 -6 653 -3
rect 302 -8 303 -6
rect 305 -8 306 -6
rect 391 -8 392 -6
rect 394 -8 395 -6
rect 560 -8 561 -6
rect 563 -8 564 -6
rect 649 -8 650 -6
rect 652 -8 653 -6
rect 212 -14 214 -12
rect 216 -14 218 -12
rect 212 -15 218 -14
rect 272 -9 297 -8
rect 203 -22 220 -18
rect 112 -44 126 -42
rect 128 -44 152 -42
rect 112 -45 152 -44
rect 168 -45 174 -41
rect 216 -27 220 -22
rect 216 -29 217 -27
rect 219 -29 220 -27
rect 125 -49 129 -45
rect 148 -49 172 -45
rect 216 -41 220 -29
rect 208 -45 220 -41
rect 208 -49 212 -45
rect 223 -49 224 -46
rect 257 -10 267 -9
rect 257 -12 263 -10
rect 265 -12 267 -10
rect 257 -13 267 -12
rect 272 -10 293 -9
rect 272 -12 273 -10
rect 275 -11 293 -10
rect 295 -11 297 -9
rect 302 -10 306 -8
rect 361 -9 386 -8
rect 275 -12 297 -11
rect 257 -17 261 -13
rect 241 -21 261 -17
rect 241 -24 245 -21
rect 239 -26 245 -24
rect 239 -28 240 -26
rect 242 -28 245 -26
rect 239 -30 245 -28
rect 241 -41 245 -30
rect 249 -26 253 -24
rect 272 -17 276 -12
rect 272 -19 273 -17
rect 275 -19 276 -17
rect 272 -21 276 -19
rect 281 -17 296 -16
rect 281 -19 283 -17
rect 285 -18 296 -17
rect 285 -19 310 -18
rect 281 -20 306 -19
rect 292 -21 306 -20
rect 308 -21 310 -19
rect 292 -22 310 -21
rect 249 -28 250 -26
rect 252 -28 253 -26
rect 249 -33 253 -28
rect 292 -33 296 -22
rect 289 -37 296 -33
rect 299 -29 303 -27
rect 299 -31 300 -29
rect 302 -31 303 -29
rect 289 -38 293 -37
rect 289 -40 290 -38
rect 292 -40 293 -38
rect 241 -42 281 -41
rect 289 -42 293 -40
rect 299 -41 303 -31
rect 241 -44 255 -42
rect 257 -44 281 -42
rect 241 -45 281 -44
rect 297 -45 303 -41
rect 25 -50 31 -49
rect 25 -52 27 -50
rect 29 -52 31 -50
rect 25 -57 31 -52
rect 36 -51 37 -49
rect 39 -51 40 -49
rect 36 -53 40 -51
rect 47 -50 53 -49
rect 47 -52 49 -50
rect 51 -52 53 -50
rect 25 -59 27 -57
rect 29 -59 31 -57
rect 47 -57 53 -52
rect 114 -50 120 -49
rect 114 -52 116 -50
rect 118 -52 120 -50
rect 47 -59 49 -57
rect 51 -59 53 -57
rect 82 -57 88 -56
rect 82 -59 84 -57
rect 86 -59 88 -57
rect 114 -57 120 -52
rect 125 -51 126 -49
rect 128 -51 129 -49
rect 125 -53 129 -51
rect 136 -50 142 -49
rect 136 -52 138 -50
rect 140 -52 142 -50
rect 114 -59 116 -57
rect 118 -59 120 -57
rect 136 -57 142 -52
rect 192 -50 212 -49
rect 192 -52 194 -50
rect 196 -52 212 -50
rect 192 -53 212 -52
rect 254 -49 258 -45
rect 277 -49 301 -45
rect 346 -10 356 -9
rect 346 -12 352 -10
rect 354 -12 356 -10
rect 346 -13 356 -12
rect 361 -10 382 -9
rect 361 -12 362 -10
rect 364 -11 382 -10
rect 384 -11 386 -9
rect 391 -10 395 -8
rect 530 -9 555 -8
rect 364 -12 386 -11
rect 346 -17 350 -13
rect 330 -21 350 -17
rect 330 -24 334 -21
rect 328 -26 334 -24
rect 328 -28 329 -26
rect 331 -28 334 -26
rect 328 -30 334 -28
rect 330 -41 334 -30
rect 338 -26 342 -24
rect 361 -17 365 -12
rect 361 -19 362 -17
rect 364 -19 365 -17
rect 361 -21 365 -19
rect 370 -17 385 -16
rect 370 -19 372 -17
rect 374 -18 385 -17
rect 374 -19 399 -18
rect 370 -20 395 -19
rect 381 -21 395 -20
rect 397 -21 399 -19
rect 381 -22 399 -21
rect 338 -28 339 -26
rect 341 -28 342 -26
rect 338 -33 342 -28
rect 381 -33 385 -22
rect 378 -37 385 -33
rect 388 -29 392 -27
rect 388 -31 389 -29
rect 391 -31 392 -29
rect 378 -38 382 -37
rect 378 -40 379 -38
rect 381 -40 382 -38
rect 330 -42 370 -41
rect 378 -42 382 -40
rect 388 -41 392 -31
rect 330 -44 344 -42
rect 346 -44 370 -42
rect 330 -45 370 -44
rect 386 -45 392 -41
rect 343 -49 347 -45
rect 366 -49 390 -45
rect 515 -10 525 -9
rect 515 -12 521 -10
rect 523 -12 525 -10
rect 515 -13 525 -12
rect 530 -10 551 -9
rect 530 -12 531 -10
rect 533 -11 551 -10
rect 553 -11 555 -9
rect 560 -10 564 -8
rect 619 -9 644 -8
rect 533 -12 555 -11
rect 515 -17 519 -13
rect 499 -21 519 -17
rect 499 -24 503 -21
rect 497 -26 503 -24
rect 497 -28 498 -26
rect 500 -28 503 -26
rect 497 -30 503 -28
rect 499 -41 503 -30
rect 507 -26 511 -24
rect 530 -17 534 -12
rect 530 -19 531 -17
rect 533 -19 534 -17
rect 530 -21 534 -19
rect 539 -17 554 -16
rect 539 -19 541 -17
rect 543 -18 554 -17
rect 543 -19 568 -18
rect 539 -20 564 -19
rect 550 -21 564 -20
rect 566 -21 568 -19
rect 550 -22 568 -21
rect 507 -28 508 -26
rect 510 -28 511 -26
rect 507 -33 511 -28
rect 550 -33 554 -22
rect 547 -37 554 -33
rect 557 -29 561 -27
rect 557 -31 558 -29
rect 560 -31 561 -29
rect 547 -38 551 -37
rect 547 -40 548 -38
rect 550 -40 551 -38
rect 499 -42 539 -41
rect 547 -42 551 -40
rect 557 -41 561 -31
rect 499 -44 513 -42
rect 515 -44 539 -42
rect 499 -45 539 -44
rect 555 -45 561 -41
rect 512 -49 516 -45
rect 535 -49 559 -45
rect 604 -10 614 -9
rect 604 -12 610 -10
rect 612 -12 614 -10
rect 604 -13 614 -12
rect 619 -10 640 -9
rect 619 -12 620 -10
rect 622 -11 640 -10
rect 642 -11 644 -9
rect 649 -10 653 -8
rect 622 -12 644 -11
rect 604 -17 608 -13
rect 588 -21 608 -17
rect 588 -24 592 -21
rect 586 -26 592 -24
rect 586 -28 587 -26
rect 589 -28 592 -26
rect 586 -30 592 -28
rect 588 -41 592 -30
rect 596 -26 600 -24
rect 619 -17 623 -12
rect 619 -19 620 -17
rect 622 -19 623 -17
rect 619 -21 623 -19
rect 628 -17 643 -16
rect 628 -19 630 -17
rect 632 -18 643 -17
rect 632 -19 657 -18
rect 628 -20 653 -19
rect 639 -21 653 -20
rect 655 -21 657 -19
rect 639 -22 657 -21
rect 596 -28 597 -26
rect 599 -28 600 -26
rect 596 -33 600 -28
rect 639 -33 643 -22
rect 636 -37 643 -33
rect 646 -29 650 -27
rect 646 -31 647 -29
rect 649 -31 650 -29
rect 636 -38 640 -37
rect 636 -40 637 -38
rect 639 -40 640 -38
rect 588 -42 628 -41
rect 636 -42 640 -40
rect 646 -41 650 -31
rect 588 -44 602 -42
rect 604 -44 628 -42
rect 588 -45 628 -44
rect 644 -45 650 -41
rect 601 -49 605 -45
rect 624 -49 648 -45
rect 243 -50 249 -49
rect 243 -52 245 -50
rect 247 -52 249 -50
rect 136 -59 138 -57
rect 140 -59 142 -57
rect 171 -57 177 -56
rect 171 -59 173 -57
rect 175 -59 177 -57
rect 210 -57 216 -56
rect 210 -59 212 -57
rect 214 -59 216 -57
rect 243 -57 249 -52
rect 254 -51 255 -49
rect 257 -51 258 -49
rect 254 -53 258 -51
rect 265 -50 271 -49
rect 265 -52 267 -50
rect 269 -52 271 -50
rect 243 -59 245 -57
rect 247 -59 249 -57
rect 265 -57 271 -52
rect 332 -50 338 -49
rect 332 -52 334 -50
rect 336 -52 338 -50
rect 265 -59 267 -57
rect 269 -59 271 -57
rect 300 -57 306 -56
rect 300 -59 302 -57
rect 304 -59 306 -57
rect 332 -57 338 -52
rect 343 -51 344 -49
rect 346 -51 347 -49
rect 343 -53 347 -51
rect 354 -50 360 -49
rect 354 -52 356 -50
rect 358 -52 360 -50
rect 332 -59 334 -57
rect 336 -59 338 -57
rect 354 -57 360 -52
rect 501 -50 507 -49
rect 501 -52 503 -50
rect 505 -52 507 -50
rect 354 -59 356 -57
rect 358 -59 360 -57
rect 389 -57 395 -56
rect 389 -59 391 -57
rect 393 -59 395 -57
rect 501 -57 507 -52
rect 512 -51 513 -49
rect 515 -51 516 -49
rect 512 -53 516 -51
rect 523 -50 529 -49
rect 523 -52 525 -50
rect 527 -52 529 -50
rect 501 -59 503 -57
rect 505 -59 507 -57
rect 523 -57 529 -52
rect 590 -50 596 -49
rect 590 -52 592 -50
rect 594 -52 596 -50
rect 523 -59 525 -57
rect 527 -59 529 -57
rect 558 -57 564 -56
rect 558 -59 560 -57
rect 562 -59 564 -57
rect 590 -57 596 -52
rect 601 -51 602 -49
rect 604 -51 605 -49
rect 601 -53 605 -51
rect 612 -50 618 -49
rect 612 -52 614 -50
rect 616 -52 618 -50
rect 590 -59 592 -57
rect 594 -59 596 -57
rect 612 -57 618 -52
rect 612 -59 614 -57
rect 616 -59 618 -57
rect 647 -57 653 -56
rect 647 -59 649 -57
rect 651 -59 653 -57
rect 18 -77 20 -75
rect 22 -77 24 -75
rect 18 -78 24 -77
rect 53 -77 55 -75
rect 57 -77 59 -75
rect 53 -82 59 -77
rect 75 -77 77 -75
rect 79 -77 81 -75
rect 53 -84 55 -82
rect 57 -84 59 -82
rect 53 -85 59 -84
rect 66 -83 70 -81
rect 66 -85 67 -83
rect 69 -85 70 -83
rect 75 -82 81 -77
rect 107 -77 109 -75
rect 111 -77 113 -75
rect 107 -78 113 -77
rect 142 -77 144 -75
rect 146 -77 148 -75
rect 75 -84 77 -82
rect 79 -84 81 -82
rect 75 -85 81 -84
rect 142 -82 148 -77
rect 164 -77 166 -75
rect 168 -77 170 -75
rect 142 -84 144 -82
rect 146 -84 148 -82
rect 142 -85 148 -84
rect 155 -83 159 -81
rect 155 -85 156 -83
rect 158 -85 159 -83
rect 164 -82 170 -77
rect 197 -77 199 -75
rect 201 -77 203 -75
rect 197 -78 203 -77
rect 236 -77 238 -75
rect 240 -77 242 -75
rect 236 -78 242 -77
rect 271 -77 273 -75
rect 275 -77 277 -75
rect 164 -84 166 -82
rect 168 -84 170 -82
rect 164 -85 170 -84
rect 23 -89 47 -85
rect 66 -89 70 -85
rect 21 -93 27 -89
rect 43 -90 83 -89
rect 43 -92 67 -90
rect 69 -92 83 -90
rect 21 -103 25 -93
rect 31 -94 35 -92
rect 43 -93 83 -92
rect 31 -96 32 -94
rect 34 -96 35 -94
rect 31 -97 35 -96
rect 21 -105 22 -103
rect 24 -105 25 -103
rect 21 -107 25 -105
rect 28 -101 35 -97
rect 28 -112 32 -101
rect 71 -106 75 -101
rect 71 -108 72 -106
rect 74 -108 75 -106
rect 14 -113 32 -112
rect 71 -110 75 -108
rect 79 -104 83 -93
rect 79 -106 85 -104
rect 79 -108 82 -106
rect 84 -108 85 -106
rect 79 -110 85 -108
rect 79 -113 83 -110
rect 14 -115 16 -113
rect 18 -114 32 -113
rect 18 -115 43 -114
rect 14 -116 39 -115
rect 28 -117 39 -116
rect 41 -117 43 -115
rect 28 -118 43 -117
rect 48 -115 52 -113
rect 48 -117 49 -115
rect 51 -117 52 -115
rect 48 -122 52 -117
rect 63 -117 83 -113
rect 63 -121 67 -117
rect 27 -123 49 -122
rect 18 -126 22 -124
rect 27 -125 29 -123
rect 31 -124 49 -123
rect 51 -124 52 -122
rect 31 -125 52 -124
rect 57 -122 67 -121
rect 57 -124 59 -122
rect 61 -124 67 -122
rect 57 -125 67 -124
rect 112 -89 136 -85
rect 155 -89 159 -85
rect 201 -82 221 -81
rect 201 -84 217 -82
rect 219 -84 221 -82
rect 201 -85 221 -84
rect 271 -82 277 -77
rect 293 -77 295 -75
rect 297 -77 299 -75
rect 271 -84 273 -82
rect 275 -84 277 -82
rect 271 -85 277 -84
rect 284 -83 288 -81
rect 284 -85 285 -83
rect 287 -85 288 -83
rect 293 -82 299 -77
rect 325 -77 327 -75
rect 329 -77 331 -75
rect 325 -78 331 -77
rect 360 -77 362 -75
rect 364 -77 366 -75
rect 293 -84 295 -82
rect 297 -84 299 -82
rect 293 -85 299 -84
rect 360 -82 366 -77
rect 382 -77 384 -75
rect 386 -77 388 -75
rect 360 -84 362 -82
rect 364 -84 366 -82
rect 360 -85 366 -84
rect 373 -83 377 -81
rect 373 -85 374 -83
rect 376 -85 377 -83
rect 382 -82 388 -77
rect 415 -77 417 -75
rect 419 -77 421 -75
rect 415 -78 421 -77
rect 454 -77 456 -75
rect 458 -77 460 -75
rect 454 -78 460 -77
rect 489 -77 491 -75
rect 493 -77 495 -75
rect 382 -84 384 -82
rect 386 -84 388 -82
rect 382 -85 388 -84
rect 110 -93 116 -89
rect 132 -90 172 -89
rect 132 -92 156 -90
rect 158 -92 172 -90
rect 110 -103 114 -93
rect 120 -94 124 -92
rect 132 -93 172 -92
rect 120 -96 121 -94
rect 123 -96 124 -94
rect 120 -97 124 -96
rect 110 -105 111 -103
rect 113 -105 114 -103
rect 110 -107 114 -105
rect 117 -101 124 -97
rect 117 -112 121 -101
rect 160 -106 164 -101
rect 160 -108 161 -106
rect 163 -108 164 -106
rect 103 -113 121 -112
rect 160 -110 164 -108
rect 168 -104 172 -93
rect 168 -106 174 -104
rect 168 -108 171 -106
rect 173 -108 174 -106
rect 168 -110 174 -108
rect 168 -113 172 -110
rect 103 -115 105 -113
rect 107 -114 121 -113
rect 107 -115 132 -114
rect 103 -116 128 -115
rect 117 -117 128 -116
rect 130 -117 132 -115
rect 117 -118 132 -117
rect 137 -115 141 -113
rect 137 -117 138 -115
rect 140 -117 141 -115
rect 137 -122 141 -117
rect 152 -117 172 -113
rect 152 -121 156 -117
rect 116 -123 138 -122
rect 27 -126 52 -125
rect 107 -126 111 -124
rect 116 -125 118 -123
rect 120 -124 138 -123
rect 140 -124 141 -122
rect 120 -125 141 -124
rect 146 -122 156 -121
rect 146 -124 148 -122
rect 150 -124 156 -122
rect 146 -125 156 -124
rect 189 -88 190 -85
rect 201 -89 205 -85
rect 193 -93 205 -89
rect 193 -105 197 -93
rect 241 -89 265 -85
rect 284 -89 288 -85
rect 193 -107 194 -105
rect 196 -107 197 -105
rect 193 -112 197 -107
rect 239 -93 245 -89
rect 261 -90 301 -89
rect 261 -92 285 -90
rect 287 -92 301 -90
rect 193 -116 210 -112
rect 116 -126 141 -125
rect 195 -120 201 -119
rect 195 -122 197 -120
rect 199 -122 201 -120
rect 18 -128 19 -126
rect 21 -128 22 -126
rect 107 -128 108 -126
rect 110 -128 111 -126
rect 18 -131 22 -128
rect 74 -129 80 -128
rect 74 -131 76 -129
rect 78 -131 80 -129
rect 107 -131 111 -128
rect 163 -129 169 -128
rect 163 -131 165 -129
rect 167 -131 169 -129
rect 195 -131 201 -122
rect 206 -120 210 -116
rect 206 -122 207 -120
rect 209 -122 210 -120
rect 206 -124 210 -122
rect 215 -120 221 -119
rect 215 -122 217 -120
rect 219 -122 221 -120
rect 215 -131 221 -122
rect 239 -103 243 -93
rect 249 -94 253 -92
rect 261 -93 301 -92
rect 249 -96 250 -94
rect 252 -96 253 -94
rect 249 -97 253 -96
rect 239 -105 240 -103
rect 242 -105 243 -103
rect 239 -107 243 -105
rect 246 -101 253 -97
rect 246 -112 250 -101
rect 289 -106 293 -101
rect 289 -108 290 -106
rect 292 -108 293 -106
rect 232 -113 250 -112
rect 289 -110 293 -108
rect 297 -104 301 -93
rect 297 -106 303 -104
rect 297 -108 300 -106
rect 302 -108 303 -106
rect 297 -110 303 -108
rect 297 -113 301 -110
rect 232 -115 234 -113
rect 236 -114 250 -113
rect 236 -115 261 -114
rect 232 -116 257 -115
rect 246 -117 257 -116
rect 259 -117 261 -115
rect 246 -118 261 -117
rect 266 -115 270 -113
rect 266 -117 267 -115
rect 269 -117 270 -115
rect 266 -122 270 -117
rect 281 -117 301 -113
rect 281 -121 285 -117
rect 245 -123 267 -122
rect 236 -126 240 -124
rect 245 -125 247 -123
rect 249 -124 267 -123
rect 269 -124 270 -122
rect 249 -125 270 -124
rect 275 -122 285 -121
rect 275 -124 277 -122
rect 279 -124 285 -122
rect 275 -125 285 -124
rect 330 -89 354 -85
rect 373 -89 377 -85
rect 419 -82 439 -81
rect 419 -84 435 -82
rect 437 -84 439 -82
rect 419 -85 439 -84
rect 489 -82 495 -77
rect 511 -77 513 -75
rect 515 -77 517 -75
rect 489 -84 491 -82
rect 493 -84 495 -82
rect 489 -85 495 -84
rect 502 -83 506 -81
rect 502 -85 503 -83
rect 505 -85 506 -83
rect 511 -82 517 -77
rect 543 -77 545 -75
rect 547 -77 549 -75
rect 543 -78 549 -77
rect 578 -77 580 -75
rect 582 -77 584 -75
rect 511 -84 513 -82
rect 515 -84 517 -82
rect 511 -85 517 -84
rect 578 -82 584 -77
rect 600 -77 602 -75
rect 604 -77 606 -75
rect 578 -84 580 -82
rect 582 -84 584 -82
rect 578 -85 584 -84
rect 591 -83 595 -81
rect 591 -85 592 -83
rect 594 -85 595 -83
rect 600 -82 606 -77
rect 633 -77 635 -75
rect 637 -77 639 -75
rect 633 -78 639 -77
rect 600 -84 602 -82
rect 604 -84 606 -82
rect 600 -85 606 -84
rect 328 -93 334 -89
rect 350 -90 390 -89
rect 350 -92 374 -90
rect 376 -92 390 -90
rect 328 -103 332 -93
rect 338 -94 342 -92
rect 350 -93 390 -92
rect 338 -96 339 -94
rect 341 -96 342 -94
rect 338 -97 342 -96
rect 328 -105 329 -103
rect 331 -105 332 -103
rect 328 -107 332 -105
rect 335 -101 342 -97
rect 335 -112 339 -101
rect 378 -106 382 -101
rect 378 -108 379 -106
rect 381 -108 382 -106
rect 321 -113 339 -112
rect 378 -110 382 -108
rect 386 -104 390 -93
rect 386 -106 392 -104
rect 386 -108 389 -106
rect 391 -108 392 -106
rect 386 -110 392 -108
rect 386 -113 390 -110
rect 321 -115 323 -113
rect 325 -114 339 -113
rect 325 -115 350 -114
rect 321 -116 346 -115
rect 335 -117 346 -116
rect 348 -117 350 -115
rect 335 -118 350 -117
rect 355 -115 359 -113
rect 355 -117 356 -115
rect 358 -117 359 -115
rect 355 -122 359 -117
rect 370 -117 390 -113
rect 370 -121 374 -117
rect 334 -123 356 -122
rect 245 -126 270 -125
rect 325 -126 329 -124
rect 334 -125 336 -123
rect 338 -124 356 -123
rect 358 -124 359 -122
rect 338 -125 359 -124
rect 364 -122 374 -121
rect 364 -124 366 -122
rect 368 -124 374 -122
rect 364 -125 374 -124
rect 407 -88 408 -85
rect 419 -89 423 -85
rect 411 -93 423 -89
rect 411 -105 415 -93
rect 459 -89 483 -85
rect 502 -89 506 -85
rect 411 -107 412 -105
rect 414 -107 415 -105
rect 411 -112 415 -107
rect 457 -93 463 -89
rect 479 -90 519 -89
rect 479 -92 503 -90
rect 505 -92 519 -90
rect 411 -116 428 -112
rect 334 -126 359 -125
rect 413 -120 419 -119
rect 413 -122 415 -120
rect 417 -122 419 -120
rect 236 -128 237 -126
rect 239 -128 240 -126
rect 325 -128 326 -126
rect 328 -128 329 -126
rect 236 -131 240 -128
rect 292 -129 298 -128
rect 292 -131 294 -129
rect 296 -131 298 -129
rect 325 -131 329 -128
rect 381 -129 387 -128
rect 381 -131 383 -129
rect 385 -131 387 -129
rect 413 -131 419 -122
rect 424 -120 428 -116
rect 424 -122 425 -120
rect 427 -122 428 -120
rect 424 -124 428 -122
rect 433 -120 439 -119
rect 433 -122 435 -120
rect 437 -122 439 -120
rect 433 -131 439 -122
rect 457 -103 461 -93
rect 467 -94 471 -92
rect 479 -93 519 -92
rect 467 -96 468 -94
rect 470 -96 471 -94
rect 467 -97 471 -96
rect 457 -105 458 -103
rect 460 -105 461 -103
rect 457 -107 461 -105
rect 464 -101 471 -97
rect 464 -112 468 -101
rect 507 -106 511 -101
rect 507 -108 508 -106
rect 510 -108 511 -106
rect 450 -113 468 -112
rect 507 -110 511 -108
rect 515 -104 519 -93
rect 515 -106 521 -104
rect 515 -108 518 -106
rect 520 -108 521 -106
rect 515 -110 521 -108
rect 515 -113 519 -110
rect 450 -115 452 -113
rect 454 -114 468 -113
rect 454 -115 479 -114
rect 450 -116 475 -115
rect 464 -117 475 -116
rect 477 -117 479 -115
rect 464 -118 479 -117
rect 484 -115 488 -113
rect 484 -117 485 -115
rect 487 -117 488 -115
rect 484 -122 488 -117
rect 499 -117 519 -113
rect 499 -121 503 -117
rect 463 -123 485 -122
rect 454 -126 458 -124
rect 463 -125 465 -123
rect 467 -124 485 -123
rect 487 -124 488 -122
rect 467 -125 488 -124
rect 493 -122 503 -121
rect 493 -124 495 -122
rect 497 -124 503 -122
rect 493 -125 503 -124
rect 548 -89 572 -85
rect 591 -89 595 -85
rect 637 -82 657 -81
rect 637 -84 653 -82
rect 655 -84 657 -82
rect 637 -85 657 -84
rect 546 -93 552 -89
rect 568 -90 608 -89
rect 568 -92 592 -90
rect 594 -92 608 -90
rect 546 -103 550 -93
rect 556 -94 560 -92
rect 568 -93 608 -92
rect 556 -96 557 -94
rect 559 -96 560 -94
rect 556 -97 560 -96
rect 546 -105 547 -103
rect 549 -105 550 -103
rect 546 -107 550 -105
rect 553 -101 560 -97
rect 553 -112 557 -101
rect 596 -106 600 -101
rect 596 -108 597 -106
rect 599 -108 600 -106
rect 539 -113 557 -112
rect 596 -110 600 -108
rect 604 -104 608 -93
rect 604 -106 610 -104
rect 604 -108 607 -106
rect 609 -108 610 -106
rect 604 -110 610 -108
rect 604 -113 608 -110
rect 539 -115 541 -113
rect 543 -114 557 -113
rect 543 -115 568 -114
rect 539 -116 564 -115
rect 553 -117 564 -116
rect 566 -117 568 -115
rect 553 -118 568 -117
rect 573 -115 577 -113
rect 573 -117 574 -115
rect 576 -117 577 -115
rect 573 -122 577 -117
rect 588 -117 608 -113
rect 588 -121 592 -117
rect 552 -123 574 -122
rect 463 -126 488 -125
rect 543 -126 547 -124
rect 552 -125 554 -123
rect 556 -124 574 -123
rect 576 -124 577 -122
rect 556 -125 577 -124
rect 582 -122 592 -121
rect 582 -124 584 -122
rect 586 -124 592 -122
rect 582 -125 592 -124
rect 625 -88 626 -85
rect 637 -89 641 -85
rect 629 -93 641 -89
rect 629 -105 633 -93
rect 629 -107 630 -105
rect 632 -107 633 -105
rect 629 -112 633 -107
rect 629 -116 646 -112
rect 552 -126 577 -125
rect 631 -120 637 -119
rect 631 -122 633 -120
rect 635 -122 637 -120
rect 454 -128 455 -126
rect 457 -128 458 -126
rect 543 -128 544 -126
rect 546 -128 547 -126
rect 454 -131 458 -128
rect 510 -129 516 -128
rect 510 -131 512 -129
rect 514 -131 516 -129
rect 543 -131 547 -128
rect 599 -129 605 -128
rect 599 -131 601 -129
rect 603 -131 605 -129
rect 631 -131 637 -122
rect 642 -120 646 -116
rect 642 -122 643 -120
rect 645 -122 646 -120
rect 642 -124 646 -122
rect 651 -120 657 -119
rect 651 -122 653 -120
rect 655 -122 657 -120
rect 651 -131 657 -122
rect 232 -156 238 -147
rect 232 -158 234 -156
rect 236 -158 238 -156
rect 232 -159 238 -158
rect 243 -156 247 -154
rect 243 -158 244 -156
rect 246 -158 247 -156
rect 243 -162 247 -158
rect 252 -156 258 -147
rect 295 -149 297 -147
rect 299 -149 301 -147
rect 295 -150 301 -149
rect 353 -150 357 -147
rect 395 -149 397 -147
rect 399 -149 401 -147
rect 395 -150 401 -149
rect 453 -150 457 -147
rect 353 -152 354 -150
rect 356 -152 357 -150
rect 453 -152 454 -150
rect 456 -152 457 -150
rect 252 -158 254 -156
rect 256 -158 258 -156
rect 252 -159 258 -158
rect 323 -153 348 -152
rect 243 -166 260 -162
rect 256 -171 260 -166
rect 256 -173 257 -171
rect 259 -173 260 -171
rect 256 -185 260 -173
rect 248 -189 260 -185
rect 248 -193 252 -189
rect 263 -193 264 -190
rect 308 -154 318 -153
rect 308 -156 314 -154
rect 316 -156 318 -154
rect 308 -157 318 -156
rect 323 -154 344 -153
rect 323 -156 324 -154
rect 326 -155 344 -154
rect 346 -155 348 -153
rect 353 -154 357 -152
rect 423 -153 448 -152
rect 326 -156 348 -155
rect 308 -161 312 -157
rect 292 -165 312 -161
rect 292 -168 296 -165
rect 290 -170 296 -168
rect 290 -172 291 -170
rect 293 -172 296 -170
rect 290 -174 296 -172
rect 292 -185 296 -174
rect 300 -170 304 -168
rect 323 -161 327 -156
rect 323 -163 324 -161
rect 326 -163 327 -161
rect 323 -165 327 -163
rect 332 -161 347 -160
rect 332 -163 334 -161
rect 336 -162 347 -161
rect 336 -163 361 -162
rect 332 -164 357 -163
rect 343 -165 357 -164
rect 359 -165 361 -163
rect 343 -166 361 -165
rect 300 -172 301 -170
rect 303 -172 304 -170
rect 300 -177 304 -172
rect 343 -177 347 -166
rect 340 -181 347 -177
rect 350 -173 354 -171
rect 350 -175 351 -173
rect 353 -175 354 -173
rect 340 -182 344 -181
rect 340 -184 341 -182
rect 343 -184 344 -182
rect 292 -186 332 -185
rect 340 -186 344 -184
rect 350 -185 354 -175
rect 292 -188 306 -186
rect 308 -188 332 -186
rect 292 -189 332 -188
rect 348 -189 354 -185
rect 232 -194 252 -193
rect 232 -196 234 -194
rect 236 -196 252 -194
rect 232 -197 252 -196
rect 305 -193 309 -189
rect 328 -193 352 -189
rect 408 -154 418 -153
rect 408 -156 414 -154
rect 416 -156 418 -154
rect 408 -157 418 -156
rect 423 -154 444 -153
rect 423 -156 424 -154
rect 426 -155 444 -154
rect 446 -155 448 -153
rect 453 -154 457 -152
rect 426 -156 448 -155
rect 408 -161 412 -157
rect 392 -165 412 -161
rect 392 -168 396 -165
rect 390 -170 396 -168
rect 390 -172 391 -170
rect 393 -172 396 -170
rect 390 -174 396 -172
rect 392 -185 396 -174
rect 400 -170 404 -168
rect 423 -161 427 -156
rect 423 -163 424 -161
rect 426 -163 427 -161
rect 423 -165 427 -163
rect 432 -161 447 -160
rect 432 -163 434 -161
rect 436 -162 447 -161
rect 436 -163 461 -162
rect 432 -164 457 -163
rect 443 -165 457 -164
rect 459 -165 461 -163
rect 443 -166 461 -165
rect 400 -172 401 -170
rect 403 -172 404 -170
rect 400 -177 404 -172
rect 443 -177 447 -166
rect 440 -181 447 -177
rect 450 -173 454 -171
rect 450 -175 451 -173
rect 453 -175 454 -173
rect 440 -182 444 -181
rect 440 -184 441 -182
rect 443 -184 444 -182
rect 392 -186 432 -185
rect 440 -186 444 -184
rect 450 -185 454 -175
rect 476 -156 482 -147
rect 476 -158 478 -156
rect 480 -158 482 -156
rect 476 -159 482 -158
rect 487 -156 491 -154
rect 487 -158 488 -156
rect 490 -158 491 -156
rect 487 -162 491 -158
rect 496 -156 502 -147
rect 539 -149 541 -147
rect 543 -149 545 -147
rect 539 -150 545 -149
rect 597 -150 601 -147
rect 639 -149 641 -147
rect 643 -149 645 -147
rect 639 -150 645 -149
rect 697 -150 701 -147
rect 597 -152 598 -150
rect 600 -152 601 -150
rect 697 -152 698 -150
rect 700 -152 701 -150
rect 496 -158 498 -156
rect 500 -158 502 -156
rect 496 -159 502 -158
rect 567 -153 592 -152
rect 487 -166 504 -162
rect 392 -188 406 -186
rect 408 -188 432 -186
rect 392 -189 432 -188
rect 448 -189 454 -185
rect 500 -171 504 -166
rect 500 -173 501 -171
rect 503 -173 504 -171
rect 405 -193 409 -189
rect 428 -193 452 -189
rect 500 -185 504 -173
rect 492 -189 504 -185
rect 492 -193 496 -189
rect 507 -193 508 -190
rect 552 -154 562 -153
rect 552 -156 558 -154
rect 560 -156 562 -154
rect 552 -157 562 -156
rect 567 -154 588 -153
rect 567 -156 568 -154
rect 570 -155 588 -154
rect 590 -155 592 -153
rect 597 -154 601 -152
rect 667 -153 692 -152
rect 570 -156 592 -155
rect 552 -161 556 -157
rect 536 -165 556 -161
rect 536 -168 540 -165
rect 534 -170 540 -168
rect 534 -172 535 -170
rect 537 -172 540 -170
rect 534 -174 540 -172
rect 536 -185 540 -174
rect 544 -170 548 -168
rect 567 -161 571 -156
rect 567 -163 568 -161
rect 570 -163 571 -161
rect 567 -165 571 -163
rect 576 -161 591 -160
rect 576 -163 578 -161
rect 580 -162 591 -161
rect 580 -163 605 -162
rect 576 -164 601 -163
rect 587 -165 601 -164
rect 603 -165 605 -163
rect 587 -166 605 -165
rect 544 -172 545 -170
rect 547 -172 548 -170
rect 544 -177 548 -172
rect 587 -177 591 -166
rect 584 -181 591 -177
rect 594 -173 598 -171
rect 594 -175 595 -173
rect 597 -175 598 -173
rect 584 -182 588 -181
rect 584 -184 585 -182
rect 587 -184 588 -182
rect 536 -186 576 -185
rect 584 -186 588 -184
rect 594 -185 598 -175
rect 536 -188 550 -186
rect 552 -188 576 -186
rect 536 -189 576 -188
rect 592 -189 598 -185
rect 294 -194 300 -193
rect 294 -196 296 -194
rect 298 -196 300 -194
rect 250 -201 256 -200
rect 250 -203 252 -201
rect 254 -203 256 -201
rect 294 -201 300 -196
rect 305 -195 306 -193
rect 308 -195 309 -193
rect 305 -197 309 -195
rect 316 -194 322 -193
rect 316 -196 318 -194
rect 320 -196 322 -194
rect 294 -203 296 -201
rect 298 -203 300 -201
rect 316 -201 322 -196
rect 394 -194 400 -193
rect 394 -196 396 -194
rect 398 -196 400 -194
rect 316 -203 318 -201
rect 320 -203 322 -201
rect 351 -201 357 -200
rect 351 -203 353 -201
rect 355 -203 357 -201
rect 394 -201 400 -196
rect 405 -195 406 -193
rect 408 -195 409 -193
rect 405 -197 409 -195
rect 416 -194 422 -193
rect 416 -196 418 -194
rect 420 -196 422 -194
rect 394 -203 396 -201
rect 398 -203 400 -201
rect 416 -201 422 -196
rect 476 -194 496 -193
rect 476 -196 478 -194
rect 480 -196 496 -194
rect 476 -197 496 -196
rect 549 -193 553 -189
rect 572 -193 596 -189
rect 652 -154 662 -153
rect 652 -156 658 -154
rect 660 -156 662 -154
rect 652 -157 662 -156
rect 667 -154 688 -153
rect 667 -156 668 -154
rect 670 -155 688 -154
rect 690 -155 692 -153
rect 697 -154 701 -152
rect 670 -156 692 -155
rect 652 -161 656 -157
rect 636 -165 656 -161
rect 636 -168 640 -165
rect 634 -170 640 -168
rect 634 -172 635 -170
rect 637 -172 640 -170
rect 634 -174 640 -172
rect 636 -185 640 -174
rect 644 -170 648 -168
rect 667 -161 671 -156
rect 667 -163 668 -161
rect 670 -163 671 -161
rect 667 -165 671 -163
rect 676 -161 691 -160
rect 676 -163 678 -161
rect 680 -162 691 -161
rect 680 -163 705 -162
rect 676 -164 701 -163
rect 687 -165 701 -164
rect 703 -165 705 -163
rect 687 -166 705 -165
rect 644 -172 645 -170
rect 647 -172 648 -170
rect 644 -177 648 -172
rect 687 -177 691 -166
rect 684 -181 691 -177
rect 694 -173 698 -171
rect 694 -175 695 -173
rect 697 -175 698 -173
rect 684 -182 688 -181
rect 684 -184 685 -182
rect 687 -184 688 -182
rect 636 -186 676 -185
rect 684 -186 688 -184
rect 694 -185 698 -175
rect 636 -188 650 -186
rect 652 -188 676 -186
rect 636 -189 676 -188
rect 692 -189 698 -185
rect 649 -193 653 -189
rect 672 -193 696 -189
rect 538 -194 544 -193
rect 538 -196 540 -194
rect 542 -196 544 -194
rect 416 -203 418 -201
rect 420 -203 422 -201
rect 451 -201 457 -200
rect 451 -203 453 -201
rect 455 -203 457 -201
rect 494 -201 500 -200
rect 494 -203 496 -201
rect 498 -203 500 -201
rect 538 -201 544 -196
rect 549 -195 550 -193
rect 552 -195 553 -193
rect 549 -197 553 -195
rect 560 -194 566 -193
rect 560 -196 562 -194
rect 564 -196 566 -194
rect 538 -203 540 -201
rect 542 -203 544 -201
rect 560 -201 566 -196
rect 638 -194 644 -193
rect 638 -196 640 -194
rect 642 -196 644 -194
rect 560 -203 562 -201
rect 564 -203 566 -201
rect 595 -201 601 -200
rect 595 -203 597 -201
rect 599 -203 601 -201
rect 638 -201 644 -196
rect 649 -195 650 -193
rect 652 -195 653 -193
rect 649 -197 653 -195
rect 660 -194 666 -193
rect 660 -196 662 -194
rect 664 -196 666 -194
rect 638 -203 640 -201
rect 642 -203 644 -201
rect 660 -201 666 -196
rect 660 -203 662 -201
rect 664 -203 666 -201
rect 695 -201 701 -200
rect 695 -203 697 -201
rect 699 -203 701 -201
rect 18 -221 20 -219
rect 22 -221 24 -219
rect 18 -222 24 -221
rect 53 -221 55 -219
rect 57 -221 59 -219
rect 53 -226 59 -221
rect 75 -221 77 -219
rect 79 -221 81 -219
rect 53 -228 55 -226
rect 57 -228 59 -226
rect 53 -229 59 -228
rect 66 -227 70 -225
rect 66 -229 67 -227
rect 69 -229 70 -227
rect 75 -226 81 -221
rect 118 -221 120 -219
rect 122 -221 124 -219
rect 118 -222 124 -221
rect 153 -221 155 -219
rect 157 -221 159 -219
rect 75 -228 77 -226
rect 79 -228 81 -226
rect 75 -229 81 -228
rect 153 -226 159 -221
rect 175 -221 177 -219
rect 179 -221 181 -219
rect 153 -228 155 -226
rect 157 -228 159 -226
rect 153 -229 159 -228
rect 166 -227 170 -225
rect 166 -229 167 -227
rect 169 -229 170 -227
rect 175 -226 181 -221
rect 219 -221 221 -219
rect 223 -221 225 -219
rect 219 -222 225 -221
rect 259 -221 261 -219
rect 263 -221 265 -219
rect 259 -222 265 -221
rect 294 -221 296 -219
rect 298 -221 300 -219
rect 175 -228 177 -226
rect 179 -228 181 -226
rect 175 -229 181 -228
rect 23 -233 47 -229
rect 66 -233 70 -229
rect 21 -237 27 -233
rect 43 -234 83 -233
rect 43 -236 67 -234
rect 69 -236 83 -234
rect 21 -247 25 -237
rect 31 -238 35 -236
rect 43 -237 83 -236
rect 31 -240 32 -238
rect 34 -240 35 -238
rect 31 -241 35 -240
rect 21 -249 22 -247
rect 24 -249 25 -247
rect 21 -251 25 -249
rect 28 -245 35 -241
rect 28 -256 32 -245
rect 71 -250 75 -245
rect 71 -252 72 -250
rect 74 -252 75 -250
rect 14 -257 32 -256
rect 71 -254 75 -252
rect 79 -248 83 -237
rect 79 -250 85 -248
rect 79 -252 82 -250
rect 84 -252 85 -250
rect 79 -254 85 -252
rect 79 -257 83 -254
rect 14 -259 16 -257
rect 18 -258 32 -257
rect 18 -259 43 -258
rect 14 -260 39 -259
rect 28 -261 39 -260
rect 41 -261 43 -259
rect 28 -262 43 -261
rect 48 -259 52 -257
rect 48 -261 49 -259
rect 51 -261 52 -259
rect 48 -266 52 -261
rect 63 -261 83 -257
rect 63 -265 67 -261
rect 27 -267 49 -266
rect 18 -270 22 -268
rect 27 -269 29 -267
rect 31 -268 49 -267
rect 51 -268 52 -266
rect 31 -269 52 -268
rect 57 -266 67 -265
rect 57 -268 59 -266
rect 61 -268 67 -266
rect 57 -269 67 -268
rect 123 -233 147 -229
rect 166 -233 170 -229
rect 223 -226 243 -225
rect 223 -228 239 -226
rect 241 -228 243 -226
rect 223 -229 243 -228
rect 294 -226 300 -221
rect 316 -221 318 -219
rect 320 -221 322 -219
rect 294 -228 296 -226
rect 298 -228 300 -226
rect 294 -229 300 -228
rect 307 -227 311 -225
rect 307 -229 308 -227
rect 310 -229 311 -227
rect 316 -226 322 -221
rect 359 -221 361 -219
rect 363 -221 365 -219
rect 359 -222 365 -221
rect 394 -221 396 -219
rect 398 -221 400 -219
rect 316 -228 318 -226
rect 320 -228 322 -226
rect 316 -229 322 -228
rect 394 -226 400 -221
rect 416 -221 418 -219
rect 420 -221 422 -219
rect 394 -228 396 -226
rect 398 -228 400 -226
rect 394 -229 400 -228
rect 407 -227 411 -225
rect 407 -229 408 -227
rect 410 -229 411 -227
rect 416 -226 422 -221
rect 460 -221 462 -219
rect 464 -221 466 -219
rect 460 -222 466 -221
rect 416 -228 418 -226
rect 420 -228 422 -226
rect 416 -229 422 -228
rect 121 -237 127 -233
rect 143 -234 183 -233
rect 143 -236 167 -234
rect 169 -236 183 -234
rect 121 -247 125 -237
rect 131 -238 135 -236
rect 143 -237 183 -236
rect 131 -240 132 -238
rect 134 -240 135 -238
rect 131 -241 135 -240
rect 121 -249 122 -247
rect 124 -249 125 -247
rect 121 -251 125 -249
rect 128 -245 135 -241
rect 128 -256 132 -245
rect 171 -250 175 -245
rect 171 -252 172 -250
rect 174 -252 175 -250
rect 114 -257 132 -256
rect 171 -254 175 -252
rect 179 -248 183 -237
rect 179 -250 185 -248
rect 179 -252 182 -250
rect 184 -252 185 -250
rect 179 -254 185 -252
rect 179 -257 183 -254
rect 114 -259 116 -257
rect 118 -258 132 -257
rect 118 -259 143 -258
rect 114 -260 139 -259
rect 128 -261 139 -260
rect 141 -261 143 -259
rect 128 -262 143 -261
rect 148 -259 152 -257
rect 148 -261 149 -259
rect 151 -261 152 -259
rect 148 -266 152 -261
rect 163 -261 183 -257
rect 163 -265 167 -261
rect 127 -267 149 -266
rect 27 -270 52 -269
rect 118 -270 122 -268
rect 127 -269 129 -267
rect 131 -268 149 -267
rect 151 -268 152 -266
rect 131 -269 152 -268
rect 157 -266 167 -265
rect 157 -268 159 -266
rect 161 -268 167 -266
rect 157 -269 167 -268
rect 211 -232 212 -229
rect 223 -233 227 -229
rect 215 -237 227 -233
rect 215 -249 219 -237
rect 264 -233 288 -229
rect 307 -233 311 -229
rect 215 -251 216 -249
rect 218 -251 219 -249
rect 215 -256 219 -251
rect 262 -237 268 -233
rect 284 -234 324 -233
rect 284 -236 308 -234
rect 310 -236 324 -234
rect 215 -260 232 -256
rect 127 -270 152 -269
rect 217 -264 223 -263
rect 217 -266 219 -264
rect 221 -266 223 -264
rect 18 -272 19 -270
rect 21 -272 22 -270
rect 118 -272 119 -270
rect 121 -272 122 -270
rect 18 -275 22 -272
rect 74 -273 80 -272
rect 74 -275 76 -273
rect 78 -275 80 -273
rect 118 -275 122 -272
rect 174 -273 180 -272
rect 174 -275 176 -273
rect 178 -275 180 -273
rect 217 -275 223 -266
rect 228 -264 232 -260
rect 228 -266 229 -264
rect 231 -266 232 -264
rect 228 -268 232 -266
rect 237 -264 243 -263
rect 237 -266 239 -264
rect 241 -266 243 -264
rect 237 -275 243 -266
rect 262 -247 266 -237
rect 272 -238 276 -236
rect 284 -237 324 -236
rect 272 -240 273 -238
rect 275 -240 276 -238
rect 272 -241 276 -240
rect 262 -249 263 -247
rect 265 -249 266 -247
rect 262 -251 266 -249
rect 269 -245 276 -241
rect 269 -256 273 -245
rect 312 -250 316 -245
rect 312 -252 313 -250
rect 315 -252 316 -250
rect 255 -257 273 -256
rect 255 -259 257 -257
rect 259 -258 273 -257
rect 259 -259 284 -258
rect 255 -260 280 -259
rect 269 -261 280 -260
rect 282 -261 284 -259
rect 269 -262 284 -261
rect 289 -259 293 -257
rect 289 -261 290 -259
rect 292 -261 293 -259
rect 289 -266 293 -261
rect 312 -254 316 -252
rect 320 -248 324 -237
rect 320 -250 326 -248
rect 320 -252 323 -250
rect 325 -252 326 -250
rect 320 -254 326 -252
rect 320 -257 324 -254
rect 304 -261 324 -257
rect 304 -265 308 -261
rect 268 -267 290 -266
rect 259 -270 263 -268
rect 268 -269 270 -267
rect 272 -268 290 -267
rect 292 -268 293 -266
rect 272 -269 293 -268
rect 298 -266 308 -265
rect 298 -268 300 -266
rect 302 -268 308 -266
rect 298 -269 308 -268
rect 364 -233 388 -229
rect 407 -233 411 -229
rect 464 -226 484 -225
rect 464 -228 480 -226
rect 482 -228 484 -226
rect 464 -229 484 -228
rect 362 -237 368 -233
rect 384 -234 424 -233
rect 384 -236 408 -234
rect 410 -236 424 -234
rect 362 -247 366 -237
rect 372 -238 376 -236
rect 384 -237 424 -236
rect 372 -240 373 -238
rect 375 -240 376 -238
rect 372 -241 376 -240
rect 362 -249 363 -247
rect 365 -249 366 -247
rect 362 -251 366 -249
rect 369 -245 376 -241
rect 369 -256 373 -245
rect 412 -250 416 -245
rect 412 -252 413 -250
rect 415 -252 416 -250
rect 355 -257 373 -256
rect 355 -259 357 -257
rect 359 -258 373 -257
rect 359 -259 384 -258
rect 355 -260 380 -259
rect 369 -261 380 -260
rect 382 -261 384 -259
rect 369 -262 384 -261
rect 389 -259 393 -257
rect 389 -261 390 -259
rect 392 -261 393 -259
rect 389 -266 393 -261
rect 412 -254 416 -252
rect 420 -248 424 -237
rect 420 -250 426 -248
rect 420 -252 423 -250
rect 425 -252 426 -250
rect 420 -254 426 -252
rect 420 -257 424 -254
rect 404 -261 424 -257
rect 404 -265 408 -261
rect 368 -267 390 -266
rect 268 -270 293 -269
rect 359 -270 363 -268
rect 368 -269 370 -267
rect 372 -268 390 -267
rect 392 -268 393 -266
rect 372 -269 393 -268
rect 398 -266 408 -265
rect 398 -268 400 -266
rect 402 -268 408 -266
rect 398 -269 408 -268
rect 452 -232 453 -229
rect 464 -233 468 -229
rect 456 -237 468 -233
rect 456 -249 460 -237
rect 456 -251 457 -249
rect 459 -251 460 -249
rect 456 -256 460 -251
rect 456 -260 473 -256
rect 368 -270 393 -269
rect 458 -264 464 -263
rect 458 -266 460 -264
rect 462 -266 464 -264
rect 259 -272 260 -270
rect 262 -272 263 -270
rect 359 -272 360 -270
rect 362 -272 363 -270
rect 259 -275 263 -272
rect 315 -273 321 -272
rect 315 -275 317 -273
rect 319 -275 321 -273
rect 359 -275 363 -272
rect 415 -273 421 -272
rect 415 -275 417 -273
rect 419 -275 421 -273
rect 458 -275 464 -266
rect 469 -264 473 -260
rect 469 -266 470 -264
rect 472 -266 473 -264
rect 469 -268 473 -266
rect 478 -264 484 -263
rect 478 -266 480 -264
rect 482 -266 484 -264
rect 478 -275 484 -266
<< via1 >>
rect 40 140 42 142
rect 84 140 86 142
rect 172 140 174 142
rect 304 140 306 142
rect 32 132 34 134
rect 120 132 122 134
rect 252 132 254 134
rect 428 132 430 134
rect 128 124 130 126
rect 216 124 218 126
rect 348 124 350 126
rect 568 124 570 126
rect 76 116 78 118
rect 208 116 210 118
rect 384 116 386 118
rect 472 116 474 118
rect 260 108 262 110
rect 392 108 394 110
rect 524 108 526 110
rect 612 108 614 110
rect 164 100 166 102
rect 340 100 342 102
rect 516 100 518 102
rect 648 100 650 102
rect 436 92 438 94
rect 480 92 482 94
rect 656 92 658 94
rect 700 92 702 94
rect 296 84 298 86
rect 560 84 562 86
rect 604 84 606 86
rect 692 84 694 86
rect -19 72 -17 74
rect 733 72 735 74
rect 32 61 34 63
rect 40 37 42 39
rect 8 29 10 31
rect 76 61 78 63
rect 84 37 86 39
rect 56 19 58 21
rect 120 61 122 63
rect 128 37 130 39
rect 97 19 99 21
rect 164 61 166 63
rect 140 36 142 38
rect 172 37 174 39
rect 208 61 210 63
rect 216 37 218 39
rect 184 27 186 29
rect 252 61 254 63
rect 228 34 230 36
rect 260 37 262 39
rect 296 61 298 63
rect 316 53 318 55
rect 304 37 306 39
rect 272 19 274 21
rect 340 61 342 63
rect 348 37 350 39
rect 384 61 386 63
rect 392 37 394 39
rect 362 19 364 21
rect 428 61 430 63
rect 436 37 438 39
rect 405 19 407 21
rect 472 61 474 63
rect 480 37 482 39
rect 448 28 450 30
rect 516 61 518 63
rect 524 37 526 39
rect 492 29 494 31
rect 560 61 562 63
rect 568 37 570 39
rect 536 28 538 30
rect 604 61 606 63
rect 612 37 614 39
rect 580 19 582 21
rect 648 61 650 63
rect 656 37 658 39
rect 629 19 631 21
rect 692 61 694 63
rect 700 37 702 39
rect -19 4 -17 6
rect 745 4 747 6
rect 48 -19 50 -17
rect 15 -34 17 -32
rect 64 -27 66 -25
rect 137 -19 139 -17
rect 106 -41 108 -39
rect 185 -20 187 -18
rect 153 -27 155 -25
rect 202 -28 204 -26
rect 201 -40 203 -38
rect 225 -36 227 -34
rect 266 -20 268 -18
rect 233 -28 235 -26
rect 282 -31 284 -29
rect 314 -26 316 -24
rect 89 -52 91 -50
rect 322 -40 324 -38
rect 346 -28 348 -26
rect 371 -27 373 -25
rect 403 -31 405 -29
rect 524 -19 526 -17
rect 492 -41 494 -39
rect 536 -36 538 -34
rect 572 -35 574 -33
rect 613 -19 615 -17
rect 581 -41 583 -39
rect 629 -27 631 -25
rect -19 -68 -17 -66
rect 732 -68 734 -66
rect 8 -105 10 -103
rect 56 -100 58 -98
rect 89 -96 91 -94
rect 56 -113 58 -111
rect 129 -105 131 -103
rect 178 -108 180 -106
rect 145 -113 147 -111
rect 97 -121 99 -119
rect 186 -116 188 -114
rect 210 -96 212 -94
rect 209 -108 211 -106
rect 226 -105 228 -103
rect 258 -100 260 -98
rect 307 -96 309 -94
rect 274 -113 276 -111
rect 347 -105 349 -103
rect 396 -108 398 -106
rect 363 -113 365 -111
rect 315 -119 317 -117
rect 404 -114 406 -112
rect 428 -96 430 -94
rect 427 -108 429 -106
rect 444 -105 446 -103
rect 484 -100 486 -98
rect 525 -96 527 -94
rect 492 -113 494 -111
rect 565 -105 567 -103
rect 614 -108 616 -106
rect 581 -113 583 -111
rect 622 -117 624 -115
rect 646 -96 648 -94
rect 645 -108 647 -106
rect -28 -136 -26 -134
rect 750 -140 752 -138
rect 242 -172 244 -170
rect 241 -184 243 -182
rect 265 -179 267 -177
rect 317 -163 319 -161
rect 284 -172 286 -170
rect 333 -175 335 -173
rect 417 -163 419 -161
rect 384 -184 386 -182
rect 434 -180 436 -178
rect 465 -175 467 -173
rect 486 -172 488 -170
rect 485 -184 487 -182
rect 561 -164 563 -162
rect 528 -172 530 -170
rect 577 -175 579 -173
rect 661 -163 663 -161
rect 628 -184 630 -182
rect 669 -180 671 -178
rect 709 -175 711 -173
rect 500 -196 502 -194
rect 737 -208 739 -206
rect -20 -212 -18 -210
rect 8 -249 10 -247
rect 67 -244 69 -242
rect 89 -240 91 -238
rect 56 -257 58 -255
rect 140 -249 142 -247
rect 189 -252 191 -250
rect 156 -257 158 -255
rect 208 -260 210 -258
rect 232 -240 234 -238
rect 231 -252 233 -250
rect 249 -249 251 -247
rect 280 -244 282 -242
rect 330 -240 332 -238
rect 297 -260 299 -258
rect 381 -249 383 -247
rect 430 -252 432 -250
rect 397 -261 399 -259
rect 473 -240 475 -238
rect 472 -252 474 -250
rect -31 -280 -29 -278
rect 719 -280 721 -278
<< via2 >>
rect -19 72 -17 74
rect 48 36 50 38
rect 153 53 155 55
rect 140 36 142 38
rect 0 29 2 31
rect -19 4 -17 6
rect -19 -68 -17 -66
rect -28 -136 -26 -134
rect -20 -212 -18 -210
rect -31 -280 -29 -278
rect 8 29 10 31
rect 64 27 66 29
rect 15 -34 17 -32
rect 89 -7 91 -5
rect 89 -96 91 -94
rect 8 -105 10 -103
rect 56 -113 58 -111
rect 137 19 139 21
rect 316 53 318 55
rect 733 72 735 74
rect 228 34 230 36
rect 380 34 382 36
rect 184 27 186 29
rect 272 19 274 21
rect 346 19 348 21
rect 274 -7 276 -5
rect 185 -20 187 -18
rect 266 -20 268 -18
rect 202 -28 204 -26
rect 233 -28 235 -26
rect 145 -34 147 -32
rect 106 -82 108 -80
rect 129 -105 131 -103
rect 97 -113 99 -111
rect 201 -40 203 -38
rect 210 -96 212 -94
rect 258 -82 260 -80
rect 225 -97 227 -95
rect 236 -97 238 -95
rect 226 -105 228 -103
rect 178 -108 180 -106
rect 209 -108 211 -106
rect 225 -113 227 -111
rect 56 -121 58 -119
rect 8 -249 10 -247
rect 97 -121 99 -119
rect 186 -121 188 -119
rect 67 -136 69 -134
rect 236 -113 238 -111
rect 282 -31 284 -29
rect 362 19 364 21
rect 371 19 373 21
rect 363 10 365 12
rect 322 -40 324 -38
rect 314 -77 316 -75
rect 307 -96 309 -94
rect 347 -105 349 -103
rect 448 28 450 30
rect 484 28 486 30
rect 492 29 494 31
rect 524 29 526 31
rect 405 19 407 21
rect 380 10 382 12
rect 403 -31 405 -29
rect 428 -96 430 -94
rect 580 19 582 21
rect 613 19 615 21
rect 745 4 747 6
rect 492 -53 494 -51
rect 553 -53 555 -51
rect 492 -85 494 -83
rect 444 -105 446 -103
rect 396 -108 398 -106
rect 427 -108 429 -106
rect 525 -96 527 -94
rect 572 -85 574 -83
rect 565 -105 567 -103
rect 553 -113 555 -111
rect 561 -113 563 -111
rect 280 -121 282 -119
rect 404 -136 406 -134
rect 280 -152 282 -150
rect 293 -152 295 -150
rect 315 -151 317 -149
rect 417 -151 419 -149
rect 225 -163 227 -161
rect 242 -172 244 -170
rect 284 -172 286 -170
rect 241 -184 243 -182
rect 156 -210 158 -208
rect 89 -240 91 -238
rect 140 -249 142 -247
rect 265 -210 267 -208
rect 280 -192 282 -190
rect 232 -240 234 -238
rect 317 -163 319 -161
rect 732 -68 734 -66
rect 661 -77 663 -75
rect 646 -96 648 -94
rect 614 -108 616 -106
rect 645 -108 647 -106
rect 622 -117 624 -115
rect 669 -117 671 -115
rect 486 -172 488 -170
rect 333 -175 335 -173
rect 528 -172 530 -170
rect 465 -175 467 -173
rect 577 -175 579 -173
rect 384 -184 386 -182
rect 293 -192 295 -190
rect 750 -140 752 -138
rect 709 -175 711 -173
rect 485 -184 487 -182
rect 628 -184 630 -182
rect 434 -196 436 -194
rect 500 -196 502 -194
rect 737 -208 739 -206
rect 330 -240 332 -238
rect 473 -240 475 -238
rect 249 -249 251 -247
rect 189 -252 191 -250
rect 381 -249 383 -247
rect 231 -252 233 -250
rect 430 -252 432 -250
rect 472 -252 474 -250
rect 208 -260 210 -258
rect 297 -260 299 -258
rect 0 -282 2 -280
rect 397 -282 399 -280
rect 719 -280 721 -278
<< via3 >>
rect -19 72 -17 74
rect 733 72 735 74
rect -19 4 -17 6
rect 745 4 747 6
rect -19 -68 -17 -66
rect 732 -68 734 -66
rect -28 -136 -26 -134
rect 750 -140 752 -138
rect -20 -212 -18 -210
rect 737 -208 739 -206
rect -31 -280 -29 -278
rect 719 -280 721 -278
<< via4 >>
rect -19 72 -17 74
rect 733 72 735 74
rect -19 4 -17 6
rect 745 4 747 6
rect -19 -68 -17 -66
rect 732 -68 734 -66
rect -28 -136 -26 -134
rect 750 -140 752 -138
rect -20 -212 -18 -210
rect 737 -208 739 -206
rect -31 -280 -29 -278
rect 719 -280 721 -278
<< via5 >>
rect -107 218 -103 222
rect 826 218 830 222
rect -55 187 -51 191
rect 772 187 776 191
rect -107 71 -103 75
rect 826 71 830 75
rect -55 4 -51 8
rect 772 4 776 8
rect -107 -69 -103 -65
rect 826 -69 830 -65
rect -55 -137 -51 -133
rect 772 -140 776 -136
rect -107 -213 -103 -209
rect 826 -209 830 -205
rect -55 -280 -51 -276
rect 772 -281 776 -277
rect -55 -333 -51 -329
rect 772 -333 776 -329
rect -107 -361 -103 -357
rect 826 -361 830 -357
<< substrateopen >>
rect 700 92 702 94
<< labels >>
rlabel alu1 25 9 25 9 6 vss
rlabel alu1 25 73 25 73 6 vdd
rlabel alu1 69 9 69 9 6 vss
rlabel alu1 69 73 69 73 6 vdd
rlabel alu1 113 9 113 9 6 vss
rlabel alu1 113 73 113 73 6 vdd
rlabel alu1 157 9 157 9 6 vss
rlabel alu1 157 73 157 73 6 vdd
rlabel alu1 245 9 245 9 6 vss
rlabel alu1 245 73 245 73 6 vdd
rlabel alu1 289 9 289 9 6 vss
rlabel alu1 289 73 289 73 6 vdd
rlabel alu1 333 9 333 9 6 vss
rlabel alu1 333 73 333 73 6 vdd
rlabel alu1 201 73 201 73 6 vdd
rlabel alu1 201 9 201 9 6 vss
rlabel alu1 377 9 377 9 6 vss
rlabel alu1 377 73 377 73 6 vdd
rlabel alu1 421 9 421 9 6 vss
rlabel alu1 421 73 421 73 6 vdd
rlabel alu1 465 9 465 9 6 vss
rlabel alu1 465 73 465 73 6 vdd
rlabel alu1 509 9 509 9 6 vss
rlabel alu1 509 73 509 73 6 vdd
rlabel alu1 553 9 553 9 6 vss
rlabel alu1 553 73 553 73 6 vdd
rlabel alu1 597 9 597 9 6 vss
rlabel alu1 597 73 597 73 6 vdd
rlabel alu1 641 9 641 9 6 vss
rlabel alu1 641 73 641 73 6 vdd
rlabel alu1 685 9 685 9 6 vss
rlabel alu1 685 73 685 73 6 vdd
rlabel alu1 692 61 692 61 1 x0
rlabel alu1 669 33 669 33 1 x0y0
rlabel alu1 648 61 648 61 1 x1
rlabel alu1 657 33 657 33 1 y0
rlabel alu1 701 33 701 33 1 y0
rlabel alu1 625 33 625 33 1 x1y0
rlabel alu1 604 61 604 61 1 x0
rlabel alu1 613 34 613 34 1 y1
rlabel alu1 581 33 581 33 1 x0y1
rlabel alu1 560 61 560 61 1 x0
rlabel alu1 569 32 569 32 1 y2
rlabel alu1 537 32 537 32 1 x0y2
rlabel alu1 516 61 516 61 1 x1
rlabel alu1 493 33 493 33 1 x1y1
rlabel alu1 472 61 472 61 1 x2
rlabel alu1 481 33 481 33 1 y0
rlabel alu1 449 34 449 34 1 x2y0
rlabel alu1 428 61 428 61 1 x3
rlabel alu1 437 33 437 33 1 y0
rlabel alu1 405 34 405 34 1 x3y0
rlabel alu1 384 61 384 61 1 x2
rlabel alu1 393 33 393 33 1 y1
rlabel alu1 340 61 340 61 1 x1
rlabel alu1 296 61 296 61 1 x0
rlabel alu1 252 61 252 61 1 x3
rlabel alu1 208 61 208 61 1 x2
rlabel alu1 217 33 217 33 1 y2
rlabel alu1 185 33 185 33 1 x2y2
rlabel alu1 164 61 164 61 1 x1
rlabel alu1 173 33 173 33 1 y3
rlabel alu1 141 33 141 33 1 x1y3
rlabel alu1 120 61 120 61 1 x3
rlabel alu1 129 33 129 33 1 y2
rlabel alu1 97 34 97 34 1 x3y2
rlabel alu1 77 61 77 61 1 x2
rlabel alu1 85 33 85 33 1 y3
rlabel alu1 53 33 53 33 1 x2y3
rlabel alu1 32 61 32 61 1 x3
rlabel alu1 41 34 41 34 1 y3
rlabel alu1 9 33 9 33 1 x3y3
rlabel alu1 706 84 706 84 7 x0
rlabel alu1 706 92 706 92 7 y0
rlabel alu1 53 1 53 1 2 vss
rlabel alu1 53 -63 53 -63 2 vdd
rlabel alu1 49 -22 49 -22 1 x1y3
rlabel alu1 142 -63 142 -63 2 vdd
rlabel alu1 142 1 142 1 2 vss
rlabel alu1 186 -27 186 -27 1 s1
rlabel alu1 105 -27 105 -27 1 c1
rlabel alu1 138 -24 138 -24 1 x0y3
rlabel alu1 360 1 360 1 2 vss
rlabel alu1 360 -63 360 -63 2 vdd
rlabel alu1 271 -63 271 -63 2 vdd
rlabel alu1 271 1 271 1 2 vss
rlabel alu1 210 1 210 1 2 vss
rlabel alu1 210 -63 210 -63 2 vdd
rlabel alu1 226 -32 226 -32 1 c4
rlabel alu1 265 -27 265 -27 1 s1
rlabel alu1 356 -23 356 -23 1 x2y1
rlabel alu1 359 -35 359 -35 1 x3y0
rlabel alu1 529 1 529 1 2 vss
rlabel alu1 529 -63 529 -63 2 vdd
rlabel alu1 492 -27 492 -27 1 c3
rlabel alu1 525 -24 525 -24 1 x1y1
rlabel alu1 526 -35 526 -35 1 x0y2
rlabel alu1 618 1 618 1 2 vss
rlabel alu1 618 -63 618 -63 2 vdd
rlabel alu1 662 -27 662 -27 1 s7
rlabel alu1 581 -27 581 -27 1 c7
rlabel alu1 614 -23 614 -23 1 x0y1
rlabel alu1 617 -35 617 -35 1 x1y0
rlabel alu1 53 -135 53 -135 6 vss
rlabel alu1 53 -71 53 -71 6 vdd
rlabel alu1 142 -71 142 -71 6 vdd
rlabel alu1 142 -135 142 -135 6 vss
rlabel alu1 203 -135 203 -135 6 vss
rlabel alu1 203 -71 203 -71 6 vdd
rlabel alu1 98 -107 98 -107 1 s6
rlabel alu1 187 -103 187 -103 1 c6
rlabel alu1 49 -99 49 -99 1 x2y3
rlabel alu1 146 -116 146 -116 1 c2
rlabel alu1 421 -71 421 -71 6 vdd
rlabel alu1 421 -135 421 -135 6 vss
rlabel alu1 360 -135 360 -135 6 vss
rlabel alu1 360 -71 360 -71 6 vdd
rlabel alu1 271 -71 271 -71 6 vdd
rlabel alu1 271 -135 271 -135 6 vss
rlabel alu1 316 -107 316 -107 1 s5
rlabel alu1 405 -101 405 -101 1 c5
rlabel alu1 273 -99 273 -99 1 c1
rlabel alu1 275 -117 275 -117 1 s2
rlabel alu1 639 -71 639 -71 6 vdd
rlabel alu1 639 -135 639 -135 6 vss
rlabel alu1 578 -135 578 -135 6 vss
rlabel alu1 578 -71 578 -71 6 vdd
rlabel alu1 489 -71 489 -71 6 vdd
rlabel alu1 489 -135 489 -135 6 vss
rlabel alu1 534 -107 534 -107 1 s8
rlabel alu1 623 -104 623 -104 1 c8
rlabel alu1 573 -27 573 -27 1 s3
rlabel alu1 493 -116 493 -116 1 s3
rlabel alu1 582 -115 582 -115 1 c7
rlabel alu1 494 -143 494 -143 2 vss
rlabel alu1 494 -207 494 -207 2 vdd
rlabel alu1 566 -207 566 -207 2 vdd
rlabel alu1 566 -143 566 -143 2 vss
rlabel alu1 666 -207 666 -207 2 vdd
rlabel alu1 666 -143 666 -143 2 vss
rlabel alu1 510 -177 510 -177 1 c9
rlabel alu1 610 -171 610 -171 1 s9
rlabel alu1 560 -171 560 -171 1 c3
rlabel alu1 662 -166 662 -166 1 s4
rlabel alu1 663 -179 663 -179 1 c8
rlabel alu1 250 -143 250 -143 2 vss
rlabel alu1 250 -207 250 -207 2 vdd
rlabel alu1 322 -207 322 -207 2 vdd
rlabel alu1 322 -143 322 -143 2 vss
rlabel alu1 422 -207 422 -207 2 vdd
rlabel alu1 422 -143 422 -143 2 vss
rlabel alu1 366 -171 366 -171 1 s10
rlabel alu1 419 -179 419 -179 1 c9
rlabel alu1 418 -168 418 -168 1 s5
rlabel alu1 318 -168 318 -168 1 c4
rlabel alu1 53 -215 53 -215 6 vdd
rlabel alu1 153 -215 153 -215 6 vdd
rlabel alu1 225 -215 225 -215 6 vdd
rlabel alu1 209 -245 209 -245 1 c11
rlabel alu1 109 -252 109 -252 1 s11
rlabel alu1 157 -260 157 -260 1 c10
rlabel alu1 57 -259 57 -259 1 s6
rlabel alu1 52 -244 52 -244 1 c5
rlabel alu1 466 -215 466 -215 6 vdd
rlabel alu1 394 -215 394 -215 6 vdd
rlabel alu1 294 -215 294 -215 6 vdd
rlabel alu1 350 -251 350 -251 1 s12
rlabel alu1 450 -247 450 -247 1 c12
rlabel alu1 298 -255 298 -255 1 c11
rlabel alu1 291 -243 291 -243 1 c6
rlabel alu1 266 -167 266 -167 1 c10
rlabel alu1 503 -99 503 -99 1 x2y0
rlabel alu1 29 -11 29 -11 1 c2
rlabel alu1 87 -51 87 -51 1 s2
rlabel alu1 154 -31 154 -31 1 x1y2
rlabel alu1 361 30 361 30 1 x2y1
rlabel alu1 349 30 349 30 1 y2
rlabel alu1 317 29 317 29 1 x1y2
rlabel alu1 305 30 305 30 1 y3
rlabel alu1 273 28 273 28 1 x0y3
rlabel alu1 261 29 261 29 1 y1
rlabel alu1 229 30 229 30 1 x3y1
rlabel alu1 315 -20 315 -20 1 s4
rlabel alu1 50 -36 50 -36 1 x2y2
rlabel alu1 525 34 525 34 1 y1
<< end >>
